// SineWave Look-Up Table Method
// Nigil

// `define ASK
// `define FSK
// `define PSK

// Timescale

`timescale 1ns / 1ps

module SineWave
(
    input CLK, RESET, rEN,
    input bit,
    output reg done,
    output reg [15:0] data_pt
    
    // Check
    
    // output [7:0] chk_count_i
    
);


// Look-Up Table
// Amplitude Max Value 16'hFFFF

reg [15:00] reg_datpt_000 = 16'h0;
reg [15:00] reg_datpt_001 = 16'h0;
reg [15:00] reg_datpt_002 = 16'h0;
reg [15:00] reg_datpt_003 = 16'h0;
reg [15:00] reg_datpt_004 = 16'h0;
reg [15:00] reg_datpt_005 = 16'h0;
reg [15:00] reg_datpt_006 = 16'h0;
reg [15:00] reg_datpt_007 = 16'h0;
reg [15:00] reg_datpt_008 = 16'h0;
reg [15:00] reg_datpt_009 = 16'h0;
reg [15:00] reg_datpt_010 = 16'h0;
reg [15:00] reg_datpt_011 = 16'h0;
reg [15:00] reg_datpt_012 = 16'h0;
reg [15:00] reg_datpt_013 = 16'h0;
reg [15:00] reg_datpt_014 = 16'h0;
reg [15:00] reg_datpt_015 = 16'h0;
reg [15:00] reg_datpt_016 = 16'h0;
reg [15:00] reg_datpt_017 = 16'h0;
reg [15:00] reg_datpt_018 = 16'h0;
reg [15:00] reg_datpt_019 = 16'h0;
reg [15:00] reg_datpt_020 = 16'h0;
reg [15:00] reg_datpt_021 = 16'h0;
reg [15:00] reg_datpt_022 = 16'h0;
reg [15:00] reg_datpt_023 = 16'h0;
reg [15:00] reg_datpt_024 = 16'h0;
reg [15:00] reg_datpt_025 = 16'h0;
reg [15:00] reg_datpt_026 = 16'h0;
reg [15:00] reg_datpt_027 = 16'h0;
reg [15:00] reg_datpt_028 = 16'h0;
reg [15:00] reg_datpt_029 = 16'h0;
reg [15:00] reg_datpt_030 = 16'h0;
reg [15:00] reg_datpt_031 = 16'h0;
reg [15:00] reg_datpt_032 = 16'h0;
reg [15:00] reg_datpt_033 = 16'h0;
reg [15:00] reg_datpt_034 = 16'h0;
reg [15:00] reg_datpt_035 = 16'h0;
reg [15:00] reg_datpt_036 = 16'h0;
reg [15:00] reg_datpt_037 = 16'h0;
reg [15:00] reg_datpt_038 = 16'h0;
reg [15:00] reg_datpt_039 = 16'h0;
reg [15:00] reg_datpt_040 = 16'h0;
reg [15:00] reg_datpt_041 = 16'h0;
reg [15:00] reg_datpt_042 = 16'h0;
reg [15:00] reg_datpt_043 = 16'h0;
reg [15:00] reg_datpt_044 = 16'h0;
reg [15:00] reg_datpt_045 = 16'h0;
reg [15:00] reg_datpt_046 = 16'h0;
reg [15:00] reg_datpt_047 = 16'h0;
reg [15:00] reg_datpt_048 = 16'h0;
reg [15:00] reg_datpt_049 = 16'h0;
reg [15:00] reg_datpt_050 = 16'h0;
reg [15:00] reg_datpt_051 = 16'h0;
reg [15:00] reg_datpt_052 = 16'h0;
reg [15:00] reg_datpt_053 = 16'h0;
reg [15:00] reg_datpt_054 = 16'h0;
reg [15:00] reg_datpt_055 = 16'h0;
reg [15:00] reg_datpt_056 = 16'h0;
reg [15:00] reg_datpt_057 = 16'h0;
reg [15:00] reg_datpt_058 = 16'h0;
reg [15:00] reg_datpt_059 = 16'h0;
reg [15:00] reg_datpt_060 = 16'h0;
reg [15:00] reg_datpt_061 = 16'h0;
reg [15:00] reg_datpt_062 = 16'h0;
reg [15:00] reg_datpt_063 = 16'h0;
reg [15:00] reg_datpt_064 = 16'h0;
reg [15:00] reg_datpt_065 = 16'h0;
reg [15:00] reg_datpt_066 = 16'h0;
reg [15:00] reg_datpt_067 = 16'h0;
reg [15:00] reg_datpt_068 = 16'h0;
reg [15:00] reg_datpt_069 = 16'h0;
reg [15:00] reg_datpt_070 = 16'h0;
reg [15:00] reg_datpt_071 = 16'h0;
reg [15:00] reg_datpt_072 = 16'h0;
reg [15:00] reg_datpt_073 = 16'h0;
reg [15:00] reg_datpt_074 = 16'h0;
reg [15:00] reg_datpt_075 = 16'h0;
reg [15:00] reg_datpt_076 = 16'h0;
reg [15:00] reg_datpt_077 = 16'h0;
reg [15:00] reg_datpt_078 = 16'h0;
reg [15:00] reg_datpt_079 = 16'h0;
reg [15:00] reg_datpt_080 = 16'h0;
reg [15:00] reg_datpt_081 = 16'h0;
reg [15:00] reg_datpt_082 = 16'h0;
reg [15:00] reg_datpt_083 = 16'h0;
reg [15:00] reg_datpt_084 = 16'h0;
reg [15:00] reg_datpt_085 = 16'h0;
reg [15:00] reg_datpt_086 = 16'h0;
reg [15:00] reg_datpt_087 = 16'h0;
reg [15:00] reg_datpt_088 = 16'h0;
reg [15:00] reg_datpt_089 = 16'h0;
reg [15:00] reg_datpt_090 = 16'h0;
reg [15:00] reg_datpt_091 = 16'h0;
reg [15:00] reg_datpt_092 = 16'h0;
reg [15:00] reg_datpt_093 = 16'h0;
reg [15:00] reg_datpt_094 = 16'h0;
reg [15:00] reg_datpt_095 = 16'h0;
reg [15:00] reg_datpt_096 = 16'h0;
reg [15:00] reg_datpt_097 = 16'h0;
reg [15:00] reg_datpt_098 = 16'h0;
reg [15:00] reg_datpt_099 = 16'h0;
reg [15:00] reg_datpt_100 = 16'h0;
reg [15:00] reg_datpt_101 = 16'h0;
reg [15:00] reg_datpt_102 = 16'h0;
reg [15:00] reg_datpt_103 = 16'h0;
reg [15:00] reg_datpt_104 = 16'h0;
reg [15:00] reg_datpt_105 = 16'h0;
reg [15:00] reg_datpt_106 = 16'h0;
reg [15:00] reg_datpt_107 = 16'h0;
reg [15:00] reg_datpt_108 = 16'h0;
reg [15:00] reg_datpt_109 = 16'h0;
reg [15:00] reg_datpt_110 = 16'h0;
reg [15:00] reg_datpt_111 = 16'h0;
reg [15:00] reg_datpt_112 = 16'h0;
reg [15:00] reg_datpt_113 = 16'h0;
reg [15:00] reg_datpt_114 = 16'h0;
reg [15:00] reg_datpt_115 = 16'h0;
reg [15:00] reg_datpt_116 = 16'h0;
reg [15:00] reg_datpt_117 = 16'h0;
reg [15:00] reg_datpt_118 = 16'h0;
reg [15:00] reg_datpt_119 = 16'h0;
reg [15:00] reg_datpt_120 = 16'h0;
reg [15:00] reg_datpt_121 = 16'h0;
reg [15:00] reg_datpt_122 = 16'h0;
reg [15:00] reg_datpt_123 = 16'h0;
reg [15:00] reg_datpt_124 = 16'h0;
reg [15:00] reg_datpt_125 = 16'h0;
reg [15:00] reg_datpt_126 = 16'h0;
reg [15:00] reg_datpt_127 = 16'h0;
reg [15:00] reg_datpt_128 = 16'h0;
reg [15:00] reg_datpt_129 = 16'h0;
reg [15:00] reg_datpt_130 = 16'h0;
reg [15:00] reg_datpt_131 = 16'h0;
reg [15:00] reg_datpt_132 = 16'h0;
reg [15:00] reg_datpt_133 = 16'h0;
reg [15:00] reg_datpt_134 = 16'h0;
reg [15:00] reg_datpt_135 = 16'h0;
reg [15:00] reg_datpt_136 = 16'h0;
reg [15:00] reg_datpt_137 = 16'h0;
reg [15:00] reg_datpt_138 = 16'h0;
reg [15:00] reg_datpt_139 = 16'h0;
reg [15:00] reg_datpt_140 = 16'h0;
reg [15:00] reg_datpt_141 = 16'h0;
reg [15:00] reg_datpt_142 = 16'h0;
reg [15:00] reg_datpt_143 = 16'h0;
reg [15:00] reg_datpt_144 = 16'h0;
reg [15:00] reg_datpt_145 = 16'h0;
reg [15:00] reg_datpt_146 = 16'h0;
reg [15:00] reg_datpt_147 = 16'h0;
reg [15:00] reg_datpt_148 = 16'h0;
reg [15:00] reg_datpt_149 = 16'h0;
reg [15:00] reg_datpt_150 = 16'h0;
reg [15:00] reg_datpt_151 = 16'h0;
reg [15:00] reg_datpt_152 = 16'h0;
reg [15:00] reg_datpt_153 = 16'h0;
reg [15:00] reg_datpt_154 = 16'h0;
reg [15:00] reg_datpt_155 = 16'h0;
reg [15:00] reg_datpt_156 = 16'h0;
reg [15:00] reg_datpt_157 = 16'h0;
reg [15:00] reg_datpt_158 = 16'h0;
reg [15:00] reg_datpt_159 = 16'h0;
reg [15:00] reg_datpt_160 = 16'h0;
reg [15:00] reg_datpt_161 = 16'h0;
reg [15:00] reg_datpt_162 = 16'h0;
reg [15:00] reg_datpt_163 = 16'h0;
reg [15:00] reg_datpt_164 = 16'h0;
reg [15:00] reg_datpt_165 = 16'h0;
reg [15:00] reg_datpt_166 = 16'h0;
reg [15:00] reg_datpt_167 = 16'h0;
reg [15:00] reg_datpt_168 = 16'h0;
reg [15:00] reg_datpt_169 = 16'h0;
reg [15:00] reg_datpt_170 = 16'h0;
reg [15:00] reg_datpt_171 = 16'h0;
reg [15:00] reg_datpt_172 = 16'h0;
reg [15:00] reg_datpt_173 = 16'h0;
reg [15:00] reg_datpt_174 = 16'h0;
reg [15:00] reg_datpt_175 = 16'h0;
reg [15:00] reg_datpt_176 = 16'h0;
reg [15:00] reg_datpt_177 = 16'h0;
reg [15:00] reg_datpt_178 = 16'h0;
reg [15:00] reg_datpt_179 = 16'h0;
reg [15:00] reg_datpt_180 = 16'h0;
reg [15:00] reg_datpt_181 = 16'h0;
reg [15:00] reg_datpt_182 = 16'h0;
reg [15:00] reg_datpt_183 = 16'h0;
reg [15:00] reg_datpt_184 = 16'h0;
reg [15:00] reg_datpt_185 = 16'h0;
reg [15:00] reg_datpt_186 = 16'h0;
reg [15:00] reg_datpt_187 = 16'h0;
reg [15:00] reg_datpt_188 = 16'h0;
reg [15:00] reg_datpt_189 = 16'h0;
reg [15:00] reg_datpt_190 = 16'h0;
reg [15:00] reg_datpt_191 = 16'h0;
reg [15:00] reg_datpt_192 = 16'h0;
reg [15:00] reg_datpt_193 = 16'h0;
reg [15:00] reg_datpt_194 = 16'h0;
reg [15:00] reg_datpt_195 = 16'h0;
reg [15:00] reg_datpt_196 = 16'h0;
reg [15:00] reg_datpt_197 = 16'h0;
reg [15:00] reg_datpt_198 = 16'h0;
reg [15:00] reg_datpt_199 = 16'h0;
reg [15:00] reg_datpt_200 = 16'h0;
reg [15:00] reg_datpt_201 = 16'h0;
reg [15:00] reg_datpt_202 = 16'h0;
reg [15:00] reg_datpt_203 = 16'h0;
reg [15:00] reg_datpt_204 = 16'h0;
reg [15:00] reg_datpt_205 = 16'h0;
reg [15:00] reg_datpt_206 = 16'h0;
reg [15:00] reg_datpt_207 = 16'h0;
reg [15:00] reg_datpt_208 = 16'h0;
reg [15:00] reg_datpt_209 = 16'h0;
reg [15:00] reg_datpt_210 = 16'h0;
reg [15:00] reg_datpt_211 = 16'h0;
reg [15:00] reg_datpt_212 = 16'h0;
reg [15:00] reg_datpt_213 = 16'h0;
reg [15:00] reg_datpt_214 = 16'h0;
reg [15:00] reg_datpt_215 = 16'h0;
reg [15:00] reg_datpt_216 = 16'h0;
reg [15:00] reg_datpt_217 = 16'h0;
reg [15:00] reg_datpt_218 = 16'h0;
reg [15:00] reg_datpt_219 = 16'h0;
reg [15:00] reg_datpt_220 = 16'h0;
reg [15:00] reg_datpt_221 = 16'h0;
reg [15:00] reg_datpt_222 = 16'h0;
reg [15:00] reg_datpt_223 = 16'h0;
reg [15:00] reg_datpt_224 = 16'h0;
reg [15:00] reg_datpt_225 = 16'h0;
reg [15:00] reg_datpt_226 = 16'h0;
reg [15:00] reg_datpt_227 = 16'h0;
reg [15:00] reg_datpt_228 = 16'h0;
reg [15:00] reg_datpt_229 = 16'h0;
reg [15:00] reg_datpt_230 = 16'h0;
reg [15:00] reg_datpt_231 = 16'h0;
reg [15:00] reg_datpt_232 = 16'h0;
reg [15:00] reg_datpt_233 = 16'h0;
reg [15:00] reg_datpt_234 = 16'h0;
reg [15:00] reg_datpt_235 = 16'h0;
reg [15:00] reg_datpt_236 = 16'h0;
reg [15:00] reg_datpt_237 = 16'h0;
reg [15:00] reg_datpt_238 = 16'h0;
reg [15:00] reg_datpt_239 = 16'h0;
reg [15:00] reg_datpt_240 = 16'h0;
reg [15:00] reg_datpt_241 = 16'h0;
reg [15:00] reg_datpt_242 = 16'h0;
reg [15:00] reg_datpt_243 = 16'h0;
reg [15:00] reg_datpt_244 = 16'h0;
reg [15:00] reg_datpt_245 = 16'h0;
reg [15:00] reg_datpt_246 = 16'h0;
reg [15:00] reg_datpt_247 = 16'h0;
reg [15:00] reg_datpt_248 = 16'h0;
reg [15:00] reg_datpt_249 = 16'h0;
reg [15:00] reg_datpt_250 = 16'h0;
reg [15:00] reg_datpt_251 = 16'h0;
reg [15:00] reg_datpt_252 = 16'h0;
reg [15:00] reg_datpt_253 = 16'h0;
reg [15:00] reg_datpt_254 = 16'h0;
reg [15:00] reg_datpt_255 = 16'h0;

reg [7:0] count_i = 8'h0;

always @(posedge CLK)
begin
    if(!RESET)                        
    begin
        data_pt <= 16'h0;
    end    
    else if(RESET && rEN)                 
    begin	                        
        if(bit == 1'b1)            
        begin 
        // Bit '1', Datapoints Common for ASK, PSK and FSK
            case (count_i)
                  0 : data_pt <= 16'h7FFF;
                  1 : data_pt <= 16'hB0FB;
                  2 : data_pt <= 16'hDA81;
                  3 : data_pt <= 16'hF640;
                  4 : data_pt <= 16'hFFFF;
                  5 : data_pt <= 16'hF640;
                  6 : data_pt <= 16'hDA81;
                  7 : data_pt <= 16'hB0FB;
                  8 : data_pt <= 16'h7FFF;
                  9 : data_pt <= 16'h4F03;
                 10 : data_pt <= 16'h257D;
                 11 : data_pt <= 16'h09BE;
                 12 : data_pt <= 16'h0000;
                 13 : data_pt <= 16'h09BE;
                 14 : data_pt <= 16'h257D;
                 15 : data_pt <= 16'h4F03;
                 16 : data_pt <= 16'h7FFF;
                 17 : data_pt <= 16'hB0FB;
                 18 : data_pt <= 16'hDA81;
                 19 : data_pt <= 16'hF640;
                 20 : data_pt <= 16'hFFFF;
                 21 : data_pt <= 16'hF640;
                 22 : data_pt <= 16'hDA81;
                 23 : data_pt <= 16'hB0FB;
                 24 : data_pt <= 16'h7FFF;
                 25 : data_pt <= 16'h4F03;
                 26 : data_pt <= 16'h257D;
                 27 : data_pt <= 16'h09BE;
                 28 : data_pt <= 16'h0000;
                 29 : data_pt <= 16'h09BE;
                 30 : data_pt <= 16'h257D;
                 31 : data_pt <= 16'h4F03;
                 32 : data_pt <= 16'h7FFF;
                 33 : data_pt <= 16'hB0FB;
                 34 : data_pt <= 16'hDA81;
                 35 : data_pt <= 16'hF640;
                 36 : data_pt <= 16'hFFFF;
                 37 : data_pt <= 16'hF640;
                 38 : data_pt <= 16'hDA81;
                 39 : data_pt <= 16'hB0FB;
                 40 : data_pt <= 16'h7FFF;
                 41 : data_pt <= 16'h4F03;
                 42 : data_pt <= 16'h257D;
                 43 : data_pt <= 16'h09BE;
                 44 : data_pt <= 16'h0000;
                 45 : data_pt <= 16'h09BE;
                 46 : data_pt <= 16'h257D;
                 47 : data_pt <= 16'h4F03;
                 48 : data_pt <= 16'h7FFF;
                 49 : data_pt <= 16'hB0FB;
                 50 : data_pt <= 16'hDA81;
                 51 : data_pt <= 16'hF640;
                 52 : data_pt <= 16'hFFFF;
                 53 : data_pt <= 16'hF640;
                 54 : data_pt <= 16'hDA81;
                 55 : data_pt <= 16'hB0FB;
                 56 : data_pt <= 16'h7FFF;
                 57 : data_pt <= 16'h4F03;
                 58 : data_pt <= 16'h257D;
                 59 : data_pt <= 16'h09BE;
                 60 : data_pt <= 16'h0000;
                 61 : data_pt <= 16'h09BE;
                 62 : data_pt <= 16'h257D;
                 63 : data_pt <= 16'h4F03;
                 64 : data_pt <= 16'h7FFF;
                 65 : data_pt <= 16'hB0FB;
                 66 : data_pt <= 16'hDA81;
                 67 : data_pt <= 16'hF640;
                 68 : data_pt <= 16'hFFFF;
                 69 : data_pt <= 16'hF640;
                 70 : data_pt <= 16'hDA81;
                 71 : data_pt <= 16'hB0FB;
                 72 : data_pt <= 16'h7FFF;
                 73 : data_pt <= 16'h4F03;
                 74 : data_pt <= 16'h257D;
                 75 : data_pt <= 16'h09BE;
                 76 : data_pt <= 16'h0000;
                 77 : data_pt <= 16'h09BE;
                 78 : data_pt <= 16'h257D;
                 79 : data_pt <= 16'h4F03;
                 80 : data_pt <= 16'h7FFF;
                 81 : data_pt <= 16'hB0FB;
                 82 : data_pt <= 16'hDA81;
                 83 : data_pt <= 16'hF640;
                 84 : data_pt <= 16'hFFFF;
                 85 : data_pt <= 16'hF640;
                 86 : data_pt <= 16'hDA81;
                 87 : data_pt <= 16'hB0FB;
                 88 : data_pt <= 16'h7FFF;
                 89 : data_pt <= 16'h4F03;
                 90 : data_pt <= 16'h257D;
                 91 : data_pt <= 16'h09BE;
                 92 : data_pt <= 16'h0000;
                 93 : data_pt <= 16'h09BE;
                 94 : data_pt <= 16'h257D;
                 95 : data_pt <= 16'h4F03;
                 96 : data_pt <= 16'h7FFF;
                 97 : data_pt <= 16'hB0FB;
                 98 : data_pt <= 16'hDA81;
                 99 : data_pt <= 16'hF640;
                100 : data_pt <= 16'hFFFF;
                101 : data_pt <= 16'hF640;
                102 : data_pt <= 16'hDA81;
                103 : data_pt <= 16'hB0FB;
                104 : data_pt <= 16'h7FFF;
                105 : data_pt <= 16'h4F03;
                106 : data_pt <= 16'h257D;
                107 : data_pt <= 16'h09BE;
                108 : data_pt <= 16'h0000;
                109 : data_pt <= 16'h09BE;
                110 : data_pt <= 16'h257D;
                111 : data_pt <= 16'h4F03;
                112 : data_pt <= 16'h7FFF;
                113 : data_pt <= 16'hB0FB;
                114 : data_pt <= 16'hDA81;
                115 : data_pt <= 16'hF640;
                116 : data_pt <= 16'hFFFF;
                117 : data_pt <= 16'hF640;
                118 : data_pt <= 16'hDA81;
                119 : data_pt <= 16'hB0FB;
                120 : data_pt <= 16'h7FFF;
                121 : data_pt <= 16'h4F03;
                122 : data_pt <= 16'h257D;
                123 : data_pt <= 16'h09BE;
                124 : data_pt <= 16'h0000;
                125 : data_pt <= 16'h09BE;
                126 : data_pt <= 16'h257D;
                127 : data_pt <= 16'h4F03;
                128 : data_pt <= 16'h7FFF;
                129 : data_pt <= 16'hB0FB;
                130 : data_pt <= 16'hDA81;
                131 : data_pt <= 16'hF640;
                132 : data_pt <= 16'hFFFF;
                133 : data_pt <= 16'hF640;
                134 : data_pt <= 16'hDA81;
                135 : data_pt <= 16'hB0FB;
                136 : data_pt <= 16'h7FFF;
                137 : data_pt <= 16'h4F03;
                138 : data_pt <= 16'h257D;
                139 : data_pt <= 16'h09BE;
                140 : data_pt <= 16'h0000;
                141 : data_pt <= 16'h09BE;
                142 : data_pt <= 16'h257D;
                143 : data_pt <= 16'h4F03;
                144 : data_pt <= 16'h7FFF;
                145 : data_pt <= 16'hB0FB;
                146 : data_pt <= 16'hDA81;
                147 : data_pt <= 16'hF640;
                148 : data_pt <= 16'hFFFF;
                149 : data_pt <= 16'hF640;
                150 : data_pt <= 16'hDA81;
                151 : data_pt <= 16'hB0FB;
                152 : data_pt <= 16'h7FFF;
                153 : data_pt <= 16'h4F03;
                154 : data_pt <= 16'h257D;
                155 : data_pt <= 16'h09BE;
                156 : data_pt <= 16'h0000;
                157 : data_pt <= 16'h09BE;
                158 : data_pt <= 16'h257D;
                159 : data_pt <= 16'h4F03;
                160 : data_pt <= 16'h7FFF;
                161 : data_pt <= 16'hB0FB;
                162 : data_pt <= 16'hDA81;
                163 : data_pt <= 16'hF640;
                164 : data_pt <= 16'hFFFF;
                165 : data_pt <= 16'hF640;
                166 : data_pt <= 16'hDA81;
                167 : data_pt <= 16'hB0FB;
                168 : data_pt <= 16'h7FFF;
                169 : data_pt <= 16'h4F03;
                170 : data_pt <= 16'h257D;
                171 : data_pt <= 16'h09BE;
                172 : data_pt <= 16'h0000;
                173 : data_pt <= 16'h09BE;
                174 : data_pt <= 16'h257D;
                175 : data_pt <= 16'h4F03;
                176 : data_pt <= 16'h7FFF;
                177 : data_pt <= 16'hB0FB;
                178 : data_pt <= 16'hDA81;
                179 : data_pt <= 16'hF640;
                180 : data_pt <= 16'hFFFF;
                181 : data_pt <= 16'hF640;
                182 : data_pt <= 16'hDA81;
                183 : data_pt <= 16'hB0FB;
                184 : data_pt <= 16'h7FFF;
                185 : data_pt <= 16'h4F03;
                186 : data_pt <= 16'h257D;
                187 : data_pt <= 16'h09BE;
                188 : data_pt <= 16'h0000;
                189 : data_pt <= 16'h09BE;
                190 : data_pt <= 16'h257D;
                191 : data_pt <= 16'h4F03;
                192 : data_pt <= 16'h7FFF;
                193 : data_pt <= 16'hB0FB;
                194 : data_pt <= 16'hDA81;
                195 : data_pt <= 16'hF640;
                196 : data_pt <= 16'hFFFF;
                197 : data_pt <= 16'hF640;
                198 : data_pt <= 16'hDA81;
                199 : data_pt <= 16'hB0FB;
                200 : data_pt <= 16'h7FFF;
                201 : data_pt <= 16'h4F03;
                202 : data_pt <= 16'h257D;
                203 : data_pt <= 16'h09BE;
                204 : data_pt <= 16'h0000;
                205 : data_pt <= 16'h09BE;
                206 : data_pt <= 16'h257D;
                207 : data_pt <= 16'h4F03;
                208 : data_pt <= 16'h7FFF;
                209 : data_pt <= 16'hB0FB;
                210 : data_pt <= 16'hDA81;
                211 : data_pt <= 16'hF640;
                212 : data_pt <= 16'hFFFF;
                213 : data_pt <= 16'hF640;
                214 : data_pt <= 16'hDA81;
                215 : data_pt <= 16'hB0FB;
                216 : data_pt <= 16'h7FFF;
                217 : data_pt <= 16'h4F03;
                218 : data_pt <= 16'h257D;
                219 : data_pt <= 16'h09BE;
                220 : data_pt <= 16'h0000;
                221 : data_pt <= 16'h09BE;
                222 : data_pt <= 16'h257D;
                223 : data_pt <= 16'h4F03;
                224 : data_pt <= 16'h7FFF;
                225 : data_pt <= 16'hB0FB;
                226 : data_pt <= 16'hDA81;
                227 : data_pt <= 16'hF640;
                228 : data_pt <= 16'hFFFF;
                229 : data_pt <= 16'hF640;
                230 : data_pt <= 16'hDA81;
                231 : data_pt <= 16'hB0FB;
                232 : data_pt <= 16'h7FFF;
                233 : data_pt <= 16'h4F03;
                234 : data_pt <= 16'h257D;
                235 : data_pt <= 16'h09BE;
                236 : data_pt <= 16'h0000;
                237 : data_pt <= 16'h09BE;
                238 : data_pt <= 16'h257D;
                239 : data_pt <= 16'h4F03;
                240 : data_pt <= 16'h7FFF;
                241 : data_pt <= 16'hB0FB;
                242 : data_pt <= 16'hDA81;
                243 : data_pt <= 16'hF640;
                244 : data_pt <= 16'hFFFF;
                245 : data_pt <= 16'hF640;
                246 : data_pt <= 16'hDA81;
                247 : data_pt <= 16'hB0FB;
                248 : data_pt <= 16'h7FFF;
                249 : data_pt <= 16'h4F03;
                250 : data_pt <= 16'h257D;
                251 : data_pt <= 16'h09BE;
                252 : data_pt <= 16'h0000;
                253 : data_pt <= 16'h09BE;
                254 : data_pt <= 16'h257D;
                255 : data_pt <= 16'h4F03;
            endcase
        end     
        else if(bit == 1'b0)
        begin
            case (count_i)          
`ifdef ASK                   
                  0 : data_pt <= 16'h3FFF;
                  1 : data_pt <= 16'h587D;
                  2 : data_pt <= 16'h6D40;
                  3 : data_pt <= 16'h7B1F;
                  4 : data_pt <= 16'h7FFF;
                  5 : data_pt <= 16'h7B1F;
                  6 : data_pt <= 16'h6D40;
                  7 : data_pt <= 16'h587D;
                  8 : data_pt <= 16'h3FFF;
                  9 : data_pt <= 16'h2781;
                 10 : data_pt <= 16'h12BE;
                 11 : data_pt <= 16'h04DF;
                 12 : data_pt <= 16'h0000;
                 13 : data_pt <= 16'h04DF;
                 14 : data_pt <= 16'h12BE;
                 15 : data_pt <= 16'h2781;
                 16 : data_pt <= 16'h3FFF;
                 17 : data_pt <= 16'h587D;
                 18 : data_pt <= 16'h6D40;
                 19 : data_pt <= 16'h7B1F;
                 20 : data_pt <= 16'h7FFF;
                 21 : data_pt <= 16'h7B1F;
                 22 : data_pt <= 16'h6D40;
                 23 : data_pt <= 16'h587D;
                 24 : data_pt <= 16'h3FFF;
                 25 : data_pt <= 16'h2781;
                 26 : data_pt <= 16'h12BE;
                 27 : data_pt <= 16'h04DF;
                 28 : data_pt <= 16'h0000;
                 29 : data_pt <= 16'h04DF;
                 30 : data_pt <= 16'h12BE;
                 31 : data_pt <= 16'h2781;
                 32 : data_pt <= 16'h3FFF;
                 33 : data_pt <= 16'h587D;
                 34 : data_pt <= 16'h6D40;
                 35 : data_pt <= 16'h7B1F;
                 36 : data_pt <= 16'h7FFF;
                 37 : data_pt <= 16'h7B1F;
                 38 : data_pt <= 16'h6D40;
                 39 : data_pt <= 16'h587D;
                 40 : data_pt <= 16'h3FFF;
                 41 : data_pt <= 16'h2781;
                 42 : data_pt <= 16'h12BE;
                 43 : data_pt <= 16'h04DF;
                 44 : data_pt <= 16'h0000;
                 45 : data_pt <= 16'h04DF;
                 46 : data_pt <= 16'h12BE;
                 47 : data_pt <= 16'h2781;
                 48 : data_pt <= 16'h3FFF;
                 49 : data_pt <= 16'h587D;
                 50 : data_pt <= 16'h6D40;
                 51 : data_pt <= 16'h7B1F;
                 52 : data_pt <= 16'h7FFF;
                 53 : data_pt <= 16'h7B1F;
                 54 : data_pt <= 16'h6D40;
                 55 : data_pt <= 16'h587D;
                 56 : data_pt <= 16'h3FFF;
                 57 : data_pt <= 16'h2781;
                 58 : data_pt <= 16'h12BE;
                 59 : data_pt <= 16'h04DF;
                 60 : data_pt <= 16'h0000;
                 61 : data_pt <= 16'h04DF;
                 62 : data_pt <= 16'h12BE;
                 63 : data_pt <= 16'h2781;
                 64 : data_pt <= 16'h3FFF;
                 65 : data_pt <= 16'h587D;
                 66 : data_pt <= 16'h6D40;
                 67 : data_pt <= 16'h7B1F;
                 68 : data_pt <= 16'h7FFF;
                 69 : data_pt <= 16'h7B1F;
                 70 : data_pt <= 16'h6D40;
                 71 : data_pt <= 16'h587D;
                 72 : data_pt <= 16'h3FFF;
                 73 : data_pt <= 16'h2781;
                 74 : data_pt <= 16'h12BE;
                 75 : data_pt <= 16'h04DF;
                 76 : data_pt <= 16'h0000;
                 77 : data_pt <= 16'h04DF;
                 78 : data_pt <= 16'h12BE;
                 79 : data_pt <= 16'h2781;
                 80 : data_pt <= 16'h3FFF;
                 81 : data_pt <= 16'h587D;
                 82 : data_pt <= 16'h6D40;
                 83 : data_pt <= 16'h7B1F;
                 84 : data_pt <= 16'h7FFF;
                 85 : data_pt <= 16'h7B1F;
                 86 : data_pt <= 16'h6D40;
                 87 : data_pt <= 16'h587D;
                 88 : data_pt <= 16'h3FFF;
                 89 : data_pt <= 16'h2781;
                 90 : data_pt <= 16'h12BE;
                 91 : data_pt <= 16'h04DF;
                 92 : data_pt <= 16'h0000;
                 93 : data_pt <= 16'h04DF;
                 94 : data_pt <= 16'h12BE;
                 95 : data_pt <= 16'h2781;
                 96 : data_pt <= 16'h3FFF;
                 97 : data_pt <= 16'h587D;
                 98 : data_pt <= 16'h6D40;
                 99 : data_pt <= 16'h7B1F;
                100 : data_pt <= 16'h7FFF;
                101 : data_pt <= 16'h7B1F;
                102 : data_pt <= 16'h6D40;
                103 : data_pt <= 16'h587D;
                104 : data_pt <= 16'h3FFF;
                105 : data_pt <= 16'h2781;
                106 : data_pt <= 16'h12BE;
                107 : data_pt <= 16'h04DF;
                108 : data_pt <= 16'h0000;
                109 : data_pt <= 16'h04DF;
                110 : data_pt <= 16'h12BE;
                111 : data_pt <= 16'h2781;
                112 : data_pt <= 16'h3FFF;
                113 : data_pt <= 16'h587D;
                114 : data_pt <= 16'h6D40;
                115 : data_pt <= 16'h7B1F;
                116 : data_pt <= 16'h7FFF;
                117 : data_pt <= 16'h7B1F;
                118 : data_pt <= 16'h6D40;
                119 : data_pt <= 16'h587D;
                120 : data_pt <= 16'h3FFF;
                121 : data_pt <= 16'h2781;
                122 : data_pt <= 16'h12BE;
                123 : data_pt <= 16'h04DF;
                124 : data_pt <= 16'h0000;
                125 : data_pt <= 16'h04DF;
                126 : data_pt <= 16'h12BE;
                127 : data_pt <= 16'h2781;
                128 : data_pt <= 16'h3FFF;
                129 : data_pt <= 16'h587D;
                130 : data_pt <= 16'h6D40;
                131 : data_pt <= 16'h7B1F;
                132 : data_pt <= 16'h7FFF;
                133 : data_pt <= 16'h7B1F;
                134 : data_pt <= 16'h6D40;
                135 : data_pt <= 16'h587D;
                136 : data_pt <= 16'h3FFF;
                137 : data_pt <= 16'h2781;
                138 : data_pt <= 16'h12BE;
                139 : data_pt <= 16'h04DF;
                140 : data_pt <= 16'h0000;
                141 : data_pt <= 16'h04DF;
                142 : data_pt <= 16'h12BE;
                143 : data_pt <= 16'h2781;
                144 : data_pt <= 16'h3FFF;
                145 : data_pt <= 16'h587D;
                146 : data_pt <= 16'h6D40;
                147 : data_pt <= 16'h7B1F;
                148 : data_pt <= 16'h7FFF;
                149 : data_pt <= 16'h7B1F;
                150 : data_pt <= 16'h6D40;
                151 : data_pt <= 16'h587D;
                152 : data_pt <= 16'h3FFF;
                153 : data_pt <= 16'h2781;
                154 : data_pt <= 16'h12BE;
                155 : data_pt <= 16'h04DF;
                156 : data_pt <= 16'h0000;
                157 : data_pt <= 16'h04DF;
                158 : data_pt <= 16'h12BE;
                159 : data_pt <= 16'h2781;
                160 : data_pt <= 16'h3FFF;
                161 : data_pt <= 16'h587D;
                162 : data_pt <= 16'h6D40;
                163 : data_pt <= 16'h7B1F;
                164 : data_pt <= 16'h7FFF;
                165 : data_pt <= 16'h7B1F;
                166 : data_pt <= 16'h6D40;
                167 : data_pt <= 16'h587D;
                168 : data_pt <= 16'h3FFF;
                169 : data_pt <= 16'h2781;
                170 : data_pt <= 16'h12BE;
                171 : data_pt <= 16'h04DF;
                172 : data_pt <= 16'h0000;
                173 : data_pt <= 16'h04DF;
                174 : data_pt <= 16'h12BE;
                175 : data_pt <= 16'h2781;
                176 : data_pt <= 16'h3FFF;
                177 : data_pt <= 16'h587D;
                178 : data_pt <= 16'h6D40;
                179 : data_pt <= 16'h7B1F;
                180 : data_pt <= 16'h7FFF;
                181 : data_pt <= 16'h7B1F;
                182 : data_pt <= 16'h6D40;
                183 : data_pt <= 16'h587D;
                184 : data_pt <= 16'h3FFF;
                185 : data_pt <= 16'h2781;
                186 : data_pt <= 16'h12BE;
                187 : data_pt <= 16'h04DF;
                188 : data_pt <= 16'h0000;
                189 : data_pt <= 16'h04DF;
                190 : data_pt <= 16'h12BE;
                191 : data_pt <= 16'h2781;
                192 : data_pt <= 16'h3FFF;
                193 : data_pt <= 16'h587D;
                194 : data_pt <= 16'h6D40;
                195 : data_pt <= 16'h7B1F;
                196 : data_pt <= 16'h7FFF;
                197 : data_pt <= 16'h7B1F;
                198 : data_pt <= 16'h6D40;
                199 : data_pt <= 16'h587D;
                200 : data_pt <= 16'h3FFF;
                201 : data_pt <= 16'h2781;
                202 : data_pt <= 16'h12BE;
                203 : data_pt <= 16'h04DF;
                204 : data_pt <= 16'h0000;
                205 : data_pt <= 16'h04DF;
                206 : data_pt <= 16'h12BE;
                207 : data_pt <= 16'h2781;
                208 : data_pt <= 16'h3FFF;
                209 : data_pt <= 16'h587D;
                210 : data_pt <= 16'h6D40;
                211 : data_pt <= 16'h7B1F;
                212 : data_pt <= 16'h7FFF;
                213 : data_pt <= 16'h7B1F;
                214 : data_pt <= 16'h6D40;
                215 : data_pt <= 16'h587D;
                216 : data_pt <= 16'h3FFF;
                217 : data_pt <= 16'h2781;
                218 : data_pt <= 16'h12BE;
                219 : data_pt <= 16'h04DF;
                220 : data_pt <= 16'h0000;
                221 : data_pt <= 16'h04DF;
                222 : data_pt <= 16'h12BE;
                223 : data_pt <= 16'h2781;
                224 : data_pt <= 16'h3FFF;
                225 : data_pt <= 16'h587D;
                226 : data_pt <= 16'h6D40;
                227 : data_pt <= 16'h7B1F;
                228 : data_pt <= 16'h7FFF;
                229 : data_pt <= 16'h7B1F;
                230 : data_pt <= 16'h6D40;
                231 : data_pt <= 16'h587D;
                232 : data_pt <= 16'h3FFF;
                233 : data_pt <= 16'h2781;
                234 : data_pt <= 16'h12BE;
                235 : data_pt <= 16'h04DF;
                236 : data_pt <= 16'h0000;
                237 : data_pt <= 16'h04DF;
                238 : data_pt <= 16'h12BE;
                239 : data_pt <= 16'h2781;
                240 : data_pt <= 16'h3FFF;
                241 : data_pt <= 16'h587D;
                242 : data_pt <= 16'h6D40;
                243 : data_pt <= 16'h7B1F;
                244 : data_pt <= 16'h7FFF;
                245 : data_pt <= 16'h7B1F;
                246 : data_pt <= 16'h6D40;
                247 : data_pt <= 16'h587D;
                248 : data_pt <= 16'h3FFF;
                249 : data_pt <= 16'h2781;
                250 : data_pt <= 16'h12BE;
                251 : data_pt <= 16'h04DF;
                252 : data_pt <= 16'h0000;
                253 : data_pt <= 16'h04DF;
                254 : data_pt <= 16'h12BE;
                255 : data_pt <= 16'h2781;          
`endif

`ifdef FSK
                  0 : data_pt <= 16'h7FFF;
                  1 : data_pt <= 16'h98F8;
                  2 : data_pt <= 16'hB0FB;
                  3 : data_pt <= 16'hC71C;
                  4 : data_pt <= 16'hDA81;
                  5 : data_pt <= 16'hEA6C;
                  6 : data_pt <= 16'hF640;
                  7 : data_pt <= 16'hFD89;
                  8 : data_pt <= 16'hFFFF;
                  9 : data_pt <= 16'hFD89;
                 10 : data_pt <= 16'hF640;
                 11 : data_pt <= 16'hEA6C;
                 12 : data_pt <= 16'hDA81;
                 13 : data_pt <= 16'hC71C;
                 14 : data_pt <= 16'hB0FB;
                 15 : data_pt <= 16'h98F8;
                 16 : data_pt <= 16'h7FFF;
                 17 : data_pt <= 16'h6706;
                 18 : data_pt <= 16'h4F03;
                 19 : data_pt <= 16'h38E2;
                 20 : data_pt <= 16'h257D;
                 21 : data_pt <= 16'h1592;
                 22 : data_pt <= 16'h09BE;
                 23 : data_pt <= 16'h0275;
                 24 : data_pt <= 16'h0000;
                 25 : data_pt <= 16'h0275;
                 26 : data_pt <= 16'h09BE;
                 27 : data_pt <= 16'h1592;
                 28 : data_pt <= 16'h257D;
                 29 : data_pt <= 16'h38E2;
                 30 : data_pt <= 16'h4F03;
                 31 : data_pt <= 16'h6706;
                 32 : data_pt <= 16'h7FFF;
                 33 : data_pt <= 16'h98F8;
                 34 : data_pt <= 16'hB0FB;
                 35 : data_pt <= 16'hC71C;
                 36 : data_pt <= 16'hDA81;
                 37 : data_pt <= 16'hEA6C;
                 38 : data_pt <= 16'hF640;
                 39 : data_pt <= 16'hFD89;
                 40 : data_pt <= 16'hFFFF;
                 41 : data_pt <= 16'hFD89;
                 42 : data_pt <= 16'hF640;
                 43 : data_pt <= 16'hEA6C;
                 44 : data_pt <= 16'hDA81;
                 45 : data_pt <= 16'hC71C;
                 46 : data_pt <= 16'hB0FB;
                 47 : data_pt <= 16'h98F8;
                 48 : data_pt <= 16'h7FFF;
                 49 : data_pt <= 16'h6706;
                 50 : data_pt <= 16'h4F03;
                 51 : data_pt <= 16'h38E2;
                 52 : data_pt <= 16'h257D;
                 53 : data_pt <= 16'h1592;
                 54 : data_pt <= 16'h09BE;
                 55 : data_pt <= 16'h0275;
                 56 : data_pt <= 16'h0000;
                 57 : data_pt <= 16'h0275;
                 58 : data_pt <= 16'h09BE;
                 59 : data_pt <= 16'h1592;
                 60 : data_pt <= 16'h257D;
                 61 : data_pt <= 16'h38E2;
                 62 : data_pt <= 16'h4F03;
                 63 : data_pt <= 16'h6706;
                 64 : data_pt <= 16'h7FFF;
                 65 : data_pt <= 16'h98F8;
                 66 : data_pt <= 16'hB0FB;
                 67 : data_pt <= 16'hC71C;
                 68 : data_pt <= 16'hDA81;
                 69 : data_pt <= 16'hEA6C;
                 70 : data_pt <= 16'hF640;
                 71 : data_pt <= 16'hFD89;
                 72 : data_pt <= 16'hFFFF;
                 73 : data_pt <= 16'hFD89;
                 74 : data_pt <= 16'hF640;
                 75 : data_pt <= 16'hEA6C;
                 76 : data_pt <= 16'hDA81;
                 77 : data_pt <= 16'hC71C;
                 78 : data_pt <= 16'hB0FB;
                 79 : data_pt <= 16'h98F8;
                 80 : data_pt <= 16'h7FFF;
                 81 : data_pt <= 16'h6706;
                 82 : data_pt <= 16'h4F03;
                 83 : data_pt <= 16'h38E2;
                 84 : data_pt <= 16'h257D;
                 85 : data_pt <= 16'h1592;
                 86 : data_pt <= 16'h09BE;
                 87 : data_pt <= 16'h0275;
                 88 : data_pt <= 16'h0000;
                 89 : data_pt <= 16'h0275;
                 90 : data_pt <= 16'h09BE;
                 91 : data_pt <= 16'h1592;
                 92 : data_pt <= 16'h257D;
                 93 : data_pt <= 16'h38E2;
                 94 : data_pt <= 16'h4F03;
                 95 : data_pt <= 16'h6706;
                 96 : data_pt <= 16'h7FFF;
                 97 : data_pt <= 16'h98F8;
                 98 : data_pt <= 16'hB0FB;
                 99 : data_pt <= 16'hC71C;
                100 : data_pt <= 16'hDA81;
                101 : data_pt <= 16'hEA6C;
                102 : data_pt <= 16'hF640;
                103 : data_pt <= 16'hFD89;
                104 : data_pt <= 16'hFFFF;
                105 : data_pt <= 16'hFD89;
                106 : data_pt <= 16'hF640;
                107 : data_pt <= 16'hEA6C;
                108 : data_pt <= 16'hDA81;
                109 : data_pt <= 16'hC71C;
                110 : data_pt <= 16'hB0FB;
                111 : data_pt <= 16'h98F8;
                112 : data_pt <= 16'h7FFF;
                113 : data_pt <= 16'h6706;
                114 : data_pt <= 16'h4F03;
                115 : data_pt <= 16'h38E2;
                116 : data_pt <= 16'h257D;
                117 : data_pt <= 16'h1592;
                118 : data_pt <= 16'h09BE;
                119 : data_pt <= 16'h0275;
                120 : data_pt <= 16'h0000;
                121 : data_pt <= 16'h0275;
                122 : data_pt <= 16'h09BE;
                123 : data_pt <= 16'h1592;
                124 : data_pt <= 16'h257D;
                125 : data_pt <= 16'h38E2;
                126 : data_pt <= 16'h4F03;
                127 : data_pt <= 16'h6706;
                128 : data_pt <= 16'h7FFF;
                129 : data_pt <= 16'h98F8;
                130 : data_pt <= 16'hB0FB;
                131 : data_pt <= 16'hC71C;
                132 : data_pt <= 16'hDA81;
                133 : data_pt <= 16'hEA6C;
                134 : data_pt <= 16'hF640;
                135 : data_pt <= 16'hFD89;
                136 : data_pt <= 16'hFFFF;
                137 : data_pt <= 16'hFD89;
                138 : data_pt <= 16'hF640;
                139 : data_pt <= 16'hEA6C;
                140 : data_pt <= 16'hDA81;
                141 : data_pt <= 16'hC71C;
                142 : data_pt <= 16'hB0FB;
                143 : data_pt <= 16'h98F8;
                144 : data_pt <= 16'h7FFF;
                145 : data_pt <= 16'h6706;
                146 : data_pt <= 16'h4F03;
                147 : data_pt <= 16'h38E2;
                148 : data_pt <= 16'h257D;
                149 : data_pt <= 16'h1592;
                150 : data_pt <= 16'h09BE;
                151 : data_pt <= 16'h0275;
                152 : data_pt <= 16'h0000;
                153 : data_pt <= 16'h0275;
                154 : data_pt <= 16'h09BE;
                155 : data_pt <= 16'h1592;
                156 : data_pt <= 16'h257D;
                157 : data_pt <= 16'h38E2;
                158 : data_pt <= 16'h4F03;
                159 : data_pt <= 16'h6706;
                160 : data_pt <= 16'h7FFF;
                161 : data_pt <= 16'h98F8;
                162 : data_pt <= 16'hB0FB;
                163 : data_pt <= 16'hC71C;
                164 : data_pt <= 16'hDA81;
                165 : data_pt <= 16'hEA6C;
                166 : data_pt <= 16'hF640;
                167 : data_pt <= 16'hFD89;
                168 : data_pt <= 16'hFFFF;
                169 : data_pt <= 16'hFD89;
                170 : data_pt <= 16'hF640;
                171 : data_pt <= 16'hEA6C;
                172 : data_pt <= 16'hDA81;
                173 : data_pt <= 16'hC71C;
                174 : data_pt <= 16'hB0FB;
                175 : data_pt <= 16'h98F8;
                176 : data_pt <= 16'h7FFF;
                177 : data_pt <= 16'h6706;
                178 : data_pt <= 16'h4F03;
                179 : data_pt <= 16'h38E2;
                180 : data_pt <= 16'h257D;
                181 : data_pt <= 16'h1592;
                182 : data_pt <= 16'h09BE;
                183 : data_pt <= 16'h0275;
                184 : data_pt <= 16'h0000;
                185 : data_pt <= 16'h0275;
                186 : data_pt <= 16'h09BE;
                187 : data_pt <= 16'h1592;
                188 : data_pt <= 16'h257D;
                189 : data_pt <= 16'h38E2;
                190 : data_pt <= 16'h4F03;
                191 : data_pt <= 16'h6706;
                192 : data_pt <= 16'h7FFF;
                193 : data_pt <= 16'h98F8;
                194 : data_pt <= 16'hB0FB;
                195 : data_pt <= 16'hC71C;
                196 : data_pt <= 16'hDA81;
                197 : data_pt <= 16'hEA6C;
                198 : data_pt <= 16'hF640;
                199 : data_pt <= 16'hFD89;
                200 : data_pt <= 16'hFFFF;
                201 : data_pt <= 16'hFD89;
                202 : data_pt <= 16'hF640;
                203 : data_pt <= 16'hEA6C;
                204 : data_pt <= 16'hDA81;
                205 : data_pt <= 16'hC71C;
                206 : data_pt <= 16'hB0FB;
                207 : data_pt <= 16'h98F8;
                208 : data_pt <= 16'h7FFF;
                209 : data_pt <= 16'h6706;
                210 : data_pt <= 16'h4F03;
                211 : data_pt <= 16'h38E2;
                212 : data_pt <= 16'h257D;
                213 : data_pt <= 16'h1592;
                214 : data_pt <= 16'h09BE;
                215 : data_pt <= 16'h0275;
                216 : data_pt <= 16'h0000;
                217 : data_pt <= 16'h0275;
                218 : data_pt <= 16'h09BE;
                219 : data_pt <= 16'h1592;
                220 : data_pt <= 16'h257D;
                221 : data_pt <= 16'h38E2;
                222 : data_pt <= 16'h4F03;
                223 : data_pt <= 16'h6706;
                224 : data_pt <= 16'h7FFF;
                225 : data_pt <= 16'h98F8;
                226 : data_pt <= 16'hB0FB;
                227 : data_pt <= 16'hC71C;
                228 : data_pt <= 16'hDA81;
                229 : data_pt <= 16'hEA6C;
                230 : data_pt <= 16'hF640;
                231 : data_pt <= 16'hFD89;
                232 : data_pt <= 16'hFFFF;
                233 : data_pt <= 16'hFD89;
                234 : data_pt <= 16'hF640;
                235 : data_pt <= 16'hEA6C;
                236 : data_pt <= 16'hDA81;
                237 : data_pt <= 16'hC71C;
                238 : data_pt <= 16'hB0FB;
                239 : data_pt <= 16'h98F8;
                240 : data_pt <= 16'h7FFF;
                241 : data_pt <= 16'h6706;
                242 : data_pt <= 16'h4F03;
                243 : data_pt <= 16'h38E2;
                244 : data_pt <= 16'h257D;
                245 : data_pt <= 16'h1592;
                246 : data_pt <= 16'h09BE;
                247 : data_pt <= 16'h0275;
                248 : data_pt <= 16'h0000;
                249 : data_pt <= 16'h0275;
                250 : data_pt <= 16'h09BE;
                251 : data_pt <= 16'h1592;
                252 : data_pt <= 16'h257D;
                253 : data_pt <= 16'h38E2;
                254 : data_pt <= 16'h4F03;
                255 : data_pt <= 16'h6706;           
`endif              
    
`ifdef PSK
                  0 : data_pt <= 16'h7FFF;
                  1 : data_pt <= 16'h4F03;
                  2 : data_pt <= 16'h257D;
                  3 : data_pt <= 16'h09BE;
                  4 : data_pt <= 16'h0000;
                  5 : data_pt <= 16'h09BE;
                  6 : data_pt <= 16'h257D;
                  7 : data_pt <= 16'h4F03;
                  8 : data_pt <= 16'h7FFF;
                  9 : data_pt <= 16'hB0FB;
                 10 : data_pt <= 16'hDA81;
                 11 : data_pt <= 16'hF640;
                 12 : data_pt <= 16'hFFFF;
                 13 : data_pt <= 16'hF640;
                 14 : data_pt <= 16'hDA81;
                 15 : data_pt <= 16'hB0FB;
                 16 : data_pt <= 16'h7FFF;
                 17 : data_pt <= 16'h4F03;
                 18 : data_pt <= 16'h257D;
                 19 : data_pt <= 16'h09BE;
                 20 : data_pt <= 16'h0000;
                 21 : data_pt <= 16'h09BE;
                 22 : data_pt <= 16'h257D;
                 23 : data_pt <= 16'h4F03;
                 24 : data_pt <= 16'h7FFF;
                 25 : data_pt <= 16'hB0FB;
                 26 : data_pt <= 16'hDA81;
                 27 : data_pt <= 16'hF640;
                 28 : data_pt <= 16'hFFFF;
                 29 : data_pt <= 16'hF640;
                 30 : data_pt <= 16'hDA81;
                 31 : data_pt <= 16'hB0FB;
                 32 : data_pt <= 16'h7FFF;
                 33 : data_pt <= 16'h4F03;
                 34 : data_pt <= 16'h257D;
                 35 : data_pt <= 16'h09BE;
                 36 : data_pt <= 16'h0000;
                 37 : data_pt <= 16'h09BE;
                 38 : data_pt <= 16'h257D;
                 39 : data_pt <= 16'h4F03;
                 40 : data_pt <= 16'h7FFF;
                 41 : data_pt <= 16'hB0FB;
                 42 : data_pt <= 16'hDA81;
                 43 : data_pt <= 16'hF640;
                 44 : data_pt <= 16'hFFFF;
                 45 : data_pt <= 16'hF640;
                 46 : data_pt <= 16'hDA81;
                 47 : data_pt <= 16'hB0FB;
                 48 : data_pt <= 16'h7FFF;
                 49 : data_pt <= 16'h4F03;
                 50 : data_pt <= 16'h257D;
                 51 : data_pt <= 16'h09BE;
                 52 : data_pt <= 16'h0000;
                 53 : data_pt <= 16'h09BE;
                 54 : data_pt <= 16'h257D;
                 55 : data_pt <= 16'h4F03;
                 56 : data_pt <= 16'h7FFF;
                 57 : data_pt <= 16'hB0FB;
                 58 : data_pt <= 16'hDA81;
                 59 : data_pt <= 16'hF640;
                 60 : data_pt <= 16'hFFFF;
                 61 : data_pt <= 16'hF640;
                 62 : data_pt <= 16'hDA81;
                 63 : data_pt <= 16'hB0FB;
                 64 : data_pt <= 16'h7FFF;
                 65 : data_pt <= 16'h4F03;
                 66 : data_pt <= 16'h257D;
                 67 : data_pt <= 16'h09BE;
                 68 : data_pt <= 16'h0000;
                 69 : data_pt <= 16'h09BE;
                 70 : data_pt <= 16'h257D;
                 71 : data_pt <= 16'h4F03;
                 72 : data_pt <= 16'h7FFF;
                 73 : data_pt <= 16'hB0FB;
                 74 : data_pt <= 16'hDA81;
                 75 : data_pt <= 16'hF640;
                 76 : data_pt <= 16'hFFFF;
                 77 : data_pt <= 16'hF640;
                 78 : data_pt <= 16'hDA81;
                 79 : data_pt <= 16'hB0FB;
                 80 : data_pt <= 16'h7FFF;
                 81 : data_pt <= 16'h4F03;
                 82 : data_pt <= 16'h257D;
                 83 : data_pt <= 16'h09BE;
                 84 : data_pt <= 16'h0000;
                 85 : data_pt <= 16'h09BE;
                 86 : data_pt <= 16'h257D;
                 87 : data_pt <= 16'h4F03;
                 88 : data_pt <= 16'h7FFF;
                 89 : data_pt <= 16'hB0FB;
                 90 : data_pt <= 16'hDA81;
                 91 : data_pt <= 16'hF640;
                 92 : data_pt <= 16'hFFFF;
                 93 : data_pt <= 16'hF640;
                 94 : data_pt <= 16'hDA81;
                 95 : data_pt <= 16'hB0FB;
                 96 : data_pt <= 16'h7FFF;
                 97 : data_pt <= 16'h4F03;
                 98 : data_pt <= 16'h257D;
                 99 : data_pt <= 16'h09BE;
                100 : data_pt <= 16'h0000;
                101 : data_pt <= 16'h09BE;
                102 : data_pt <= 16'h257D;
                103 : data_pt <= 16'h4F03;
                104 : data_pt <= 16'h7FFF;
                105 : data_pt <= 16'hB0FB;
                106 : data_pt <= 16'hDA81;
                107 : data_pt <= 16'hF640;
                108 : data_pt <= 16'hFFFF;
                109 : data_pt <= 16'hF640;
                110 : data_pt <= 16'hDA81;
                111 : data_pt <= 16'hB0FB;
                112 : data_pt <= 16'h7FFF;
                113 : data_pt <= 16'h4F03;
                114 : data_pt <= 16'h257D;
                115 : data_pt <= 16'h09BE;
                116 : data_pt <= 16'h0000;
                117 : data_pt <= 16'h09BE;
                118 : data_pt <= 16'h257D;
                119 : data_pt <= 16'h4F03;
                120 : data_pt <= 16'h7FFF;
                121 : data_pt <= 16'hB0FB;
                122 : data_pt <= 16'hDA81;
                123 : data_pt <= 16'hF640;
                124 : data_pt <= 16'hFFFF;
                125 : data_pt <= 16'hF640;
                126 : data_pt <= 16'hDA81;
                127 : data_pt <= 16'hB0FB;
                128 : data_pt <= 16'h7FFF;
                129 : data_pt <= 16'h4F03;
                130 : data_pt <= 16'h257D;
                131 : data_pt <= 16'h09BE;
                132 : data_pt <= 16'h0000;
                133 : data_pt <= 16'h09BE;
                134 : data_pt <= 16'h257D;
                135 : data_pt <= 16'h4F03;
                136 : data_pt <= 16'h7FFF;
                137 : data_pt <= 16'hB0FB;
                138 : data_pt <= 16'hDA81;
                139 : data_pt <= 16'hF640;
                140 : data_pt <= 16'hFFFF;
                141 : data_pt <= 16'hF640;
                142 : data_pt <= 16'hDA81;
                143 : data_pt <= 16'hB0FB;
                144 : data_pt <= 16'h7FFF;
                145 : data_pt <= 16'h4F03;
                146 : data_pt <= 16'h257D;
                147 : data_pt <= 16'h09BE;
                148 : data_pt <= 16'h0000;
                149 : data_pt <= 16'h09BE;
                150 : data_pt <= 16'h257D;
                151 : data_pt <= 16'h4F03;
                152 : data_pt <= 16'h7FFF;
                153 : data_pt <= 16'hB0FB;
                154 : data_pt <= 16'hDA81;
                155 : data_pt <= 16'hF640;
                156 : data_pt <= 16'hFFFF;
                157 : data_pt <= 16'hF640;
                158 : data_pt <= 16'hDA81;
                159 : data_pt <= 16'hB0FB;
                160 : data_pt <= 16'h7FFF;
                161 : data_pt <= 16'h4F03;
                162 : data_pt <= 16'h257D;
                163 : data_pt <= 16'h09BE;
                164 : data_pt <= 16'h0000;
                165 : data_pt <= 16'h09BE;
                166 : data_pt <= 16'h257D;
                167 : data_pt <= 16'h4F03;
                168 : data_pt <= 16'h7FFF;
                169 : data_pt <= 16'hB0FB;
                170 : data_pt <= 16'hDA81;
                171 : data_pt <= 16'hF640;
                172 : data_pt <= 16'hFFFF;
                173 : data_pt <= 16'hF640;
                174 : data_pt <= 16'hDA81;
                175 : data_pt <= 16'hB0FB;
                176 : data_pt <= 16'h7FFF;
                177 : data_pt <= 16'h4F03;
                178 : data_pt <= 16'h257D;
                179 : data_pt <= 16'h09BE;
                180 : data_pt <= 16'h0000;
                181 : data_pt <= 16'h09BE;
                182 : data_pt <= 16'h257D;
                183 : data_pt <= 16'h4F03;
                184 : data_pt <= 16'h7FFF;
                185 : data_pt <= 16'hB0FB;
                186 : data_pt <= 16'hDA81;
                187 : data_pt <= 16'hF640;
                188 : data_pt <= 16'hFFFF;
                189 : data_pt <= 16'hF640;
                190 : data_pt <= 16'hDA81;
                191 : data_pt <= 16'hB0FB;
                192 : data_pt <= 16'h7FFF;
                193 : data_pt <= 16'h4F03;
                194 : data_pt <= 16'h257D;
                195 : data_pt <= 16'h09BE;
                196 : data_pt <= 16'h0000;
                197 : data_pt <= 16'h09BE;
                198 : data_pt <= 16'h257D;
                199 : data_pt <= 16'h4F03;
                200 : data_pt <= 16'h7FFF;
                201 : data_pt <= 16'hB0FB;
                202 : data_pt <= 16'hDA81;
                203 : data_pt <= 16'hF640;
                204 : data_pt <= 16'hFFFF;
                205 : data_pt <= 16'hF640;
                206 : data_pt <= 16'hDA81;
                207 : data_pt <= 16'hB0FB;
                208 : data_pt <= 16'h7FFF;
                209 : data_pt <= 16'h4F03;
                210 : data_pt <= 16'h257D;
                211 : data_pt <= 16'h09BE;
                212 : data_pt <= 16'h0000;
                213 : data_pt <= 16'h09BE;
                214 : data_pt <= 16'h257D;
                215 : data_pt <= 16'h4F03;
                216 : data_pt <= 16'h7FFF;
                217 : data_pt <= 16'hB0FB;
                218 : data_pt <= 16'hDA81;
                219 : data_pt <= 16'hF640;
                220 : data_pt <= 16'hFFFF;
                221 : data_pt <= 16'hF640;
                222 : data_pt <= 16'hDA81;
                223 : data_pt <= 16'hB0FB;
                224 : data_pt <= 16'h7FFF;
                225 : data_pt <= 16'h4F03;
                226 : data_pt <= 16'h257D;
                227 : data_pt <= 16'h09BE;
                228 : data_pt <= 16'h0000;
                229 : data_pt <= 16'h09BE;
                230 : data_pt <= 16'h257D;
                231 : data_pt <= 16'h4F03;
                232 : data_pt <= 16'h7FFF;
                233 : data_pt <= 16'hB0FB;
                234 : data_pt <= 16'hDA81;
                235 : data_pt <= 16'hF640;
                236 : data_pt <= 16'hFFFF;
                237 : data_pt <= 16'hF640;
                238 : data_pt <= 16'hDA81;
                239 : data_pt <= 16'hB0FB;
                240 : data_pt <= 16'h7FFF;
                241 : data_pt <= 16'h4F03;
                242 : data_pt <= 16'h257D;
                243 : data_pt <= 16'h09BE;
                244 : data_pt <= 16'h0000;
                245 : data_pt <= 16'h09BE;
                246 : data_pt <= 16'h257D;
                247 : data_pt <= 16'h4F03;
                248 : data_pt <= 16'h7FFF;
                249 : data_pt <= 16'hB0FB;
                250 : data_pt <= 16'hDA81;
                251 : data_pt <= 16'hF640;
                252 : data_pt <= 16'hFFFF;
                253 : data_pt <= 16'hF640;
                254 : data_pt <= 16'hDA81;
                255 : data_pt <= 16'hB0FB;
`endif             
            endcase         
        end
        if(count_i != 255 && RESET) begin
            done    <= 0;
            count_i <= count_i + 8'h1;  
        end
        else if(count_i == 255 && RESET) begin
            done    <= 1;
            count_i <= 0;
        end              
    end
end 


// assign chk_count_i = count_i; 

endmodule
