// SineWave for Amplitude Shift Keying (ASK)
// Nigil

// Timescale

`timescale 1ns / 1ps

module SineWave
(
    input CLK, RST,
    input Bit,
    output reg dFLAG,
    output reg [15:0] data_pt
);


// Registers - Look-Up Table
// Amplitude Max Value 16'hFFFF

reg [15:00] reg_datpt_000 = 16'h7FFF;
reg [15:00] reg_datpt_001 = 16'hB0FB;
reg [15:00] reg_datpt_002 = 16'hDA81;
reg [15:00] reg_datpt_003 = 16'hF640;
reg [15:00] reg_datpt_004 = 16'hFFFF;
reg [15:00] reg_datpt_005 = 16'hF640;
reg [15:00] reg_datpt_006 = 16'hDA81;
reg [15:00] reg_datpt_007 = 16'hB0FB;
reg [15:00] reg_datpt_008 = 16'h7FFF;
reg [15:00] reg_datpt_009 = 16'h4F03;
reg [15:00] reg_datpt_010 = 16'h257D;
reg [15:00] reg_datpt_011 = 16'h09BE;
reg [15:00] reg_datpt_012 = 16'h0000;
reg [15:00] reg_datpt_013 = 16'h09BE;
reg [15:00] reg_datpt_014 = 16'h257D;
reg [15:00] reg_datpt_015 = 16'h4F03;
reg [15:00] reg_datpt_016 = 16'h7FFF;
reg [15:00] reg_datpt_017 = 16'hB0FB;
reg [15:00] reg_datpt_018 = 16'hDA81;
reg [15:00] reg_datpt_019 = 16'hF640;
reg [15:00] reg_datpt_020 = 16'hFFFF;
reg [15:00] reg_datpt_021 = 16'hF640;
reg [15:00] reg_datpt_022 = 16'hDA81;
reg [15:00] reg_datpt_023 = 16'hB0FB;
reg [15:00] reg_datpt_024 = 16'h7FFF;
reg [15:00] reg_datpt_025 = 16'h4F03;
reg [15:00] reg_datpt_026 = 16'h257D;
reg [15:00] reg_datpt_027 = 16'h09BE;
reg [15:00] reg_datpt_028 = 16'h0000;
reg [15:00] reg_datpt_029 = 16'h09BE;
reg [15:00] reg_datpt_030 = 16'h257D;
reg [15:00] reg_datpt_031 = 16'h4F03;
reg [15:00] reg_datpt_032 = 16'h7FFF;
reg [15:00] reg_datpt_033 = 16'hB0FB;
reg [15:00] reg_datpt_034 = 16'hDA81;
reg [15:00] reg_datpt_035 = 16'hF640;
reg [15:00] reg_datpt_036 = 16'hFFFF;
reg [15:00] reg_datpt_037 = 16'hF640;
reg [15:00] reg_datpt_038 = 16'hDA81;
reg [15:00] reg_datpt_039 = 16'hB0FB;
reg [15:00] reg_datpt_040 = 16'h7FFF;
reg [15:00] reg_datpt_041 = 16'h4F03;
reg [15:00] reg_datpt_042 = 16'h257D;
reg [15:00] reg_datpt_043 = 16'h09BE;
reg [15:00] reg_datpt_044 = 16'h0000;
reg [15:00] reg_datpt_045 = 16'h09BE;
reg [15:00] reg_datpt_046 = 16'h257D;
reg [15:00] reg_datpt_047 = 16'h4F03;
reg [15:00] reg_datpt_048 = 16'h7FFF;
reg [15:00] reg_datpt_049 = 16'hB0FB;
reg [15:00] reg_datpt_050 = 16'hDA81;
reg [15:00] reg_datpt_051 = 16'hF640;
reg [15:00] reg_datpt_052 = 16'hFFFF;
reg [15:00] reg_datpt_053 = 16'hF640;
reg [15:00] reg_datpt_054 = 16'hDA81;
reg [15:00] reg_datpt_055 = 16'hB0FB;
reg [15:00] reg_datpt_056 = 16'h7FFF;
reg [15:00] reg_datpt_057 = 16'h4F03;
reg [15:00] reg_datpt_058 = 16'h257D;
reg [15:00] reg_datpt_059 = 16'h09BE;
reg [15:00] reg_datpt_060 = 16'h0000;
reg [15:00] reg_datpt_061 = 16'h09BE;
reg [15:00] reg_datpt_062 = 16'h257D;
reg [15:00] reg_datpt_063 = 16'h4F03;
reg [15:00] reg_datpt_064 = 16'h7FFF;
reg [15:00] reg_datpt_065 = 16'hB0FB;
reg [15:00] reg_datpt_066 = 16'hDA81;
reg [15:00] reg_datpt_067 = 16'hF640;
reg [15:00] reg_datpt_068 = 16'hFFFF;
reg [15:00] reg_datpt_069 = 16'hF640;
reg [15:00] reg_datpt_070 = 16'hDA81;
reg [15:00] reg_datpt_071 = 16'hB0FB;
reg [15:00] reg_datpt_072 = 16'h7FFF;
reg [15:00] reg_datpt_073 = 16'h4F03;
reg [15:00] reg_datpt_074 = 16'h257D;
reg [15:00] reg_datpt_075 = 16'h09BE;
reg [15:00] reg_datpt_076 = 16'h0000;
reg [15:00] reg_datpt_077 = 16'h09BE;
reg [15:00] reg_datpt_078 = 16'h257D;
reg [15:00] reg_datpt_079 = 16'h4F03;
reg [15:00] reg_datpt_080 = 16'h7FFF;
reg [15:00] reg_datpt_081 = 16'hB0FB;
reg [15:00] reg_datpt_082 = 16'hDA81;
reg [15:00] reg_datpt_083 = 16'hF640;
reg [15:00] reg_datpt_084 = 16'hFFFF;
reg [15:00] reg_datpt_085 = 16'hF640;
reg [15:00] reg_datpt_086 = 16'hDA81;
reg [15:00] reg_datpt_087 = 16'hB0FB;
reg [15:00] reg_datpt_088 = 16'h7FFF;
reg [15:00] reg_datpt_089 = 16'h4F03;
reg [15:00] reg_datpt_090 = 16'h257D;
reg [15:00] reg_datpt_091 = 16'h09BE;
reg [15:00] reg_datpt_092 = 16'h0000;
reg [15:00] reg_datpt_093 = 16'h09BE;
reg [15:00] reg_datpt_094 = 16'h257D;
reg [15:00] reg_datpt_095 = 16'h4F03;
reg [15:00] reg_datpt_096 = 16'h7FFF;
reg [15:00] reg_datpt_097 = 16'hB0FB;
reg [15:00] reg_datpt_098 = 16'hDA81;
reg [15:00] reg_datpt_099 = 16'hF640;
reg [15:00] reg_datpt_100 = 16'hFFFF;
reg [15:00] reg_datpt_101 = 16'hF640;
reg [15:00] reg_datpt_102 = 16'hDA81;
reg [15:00] reg_datpt_103 = 16'hB0FB;
reg [15:00] reg_datpt_104 = 16'h7FFF;
reg [15:00] reg_datpt_105 = 16'h4F03;
reg [15:00] reg_datpt_106 = 16'h257D;
reg [15:00] reg_datpt_107 = 16'h09BE;
reg [15:00] reg_datpt_108 = 16'h0000;
reg [15:00] reg_datpt_109 = 16'h09BE;
reg [15:00] reg_datpt_110 = 16'h257D;
reg [15:00] reg_datpt_111 = 16'h4F03;
reg [15:00] reg_datpt_112 = 16'h7FFF;
reg [15:00] reg_datpt_113 = 16'hB0FB;
reg [15:00] reg_datpt_114 = 16'hDA81;
reg [15:00] reg_datpt_115 = 16'hF640;
reg [15:00] reg_datpt_116 = 16'hFFFF;
reg [15:00] reg_datpt_117 = 16'hF640;
reg [15:00] reg_datpt_118 = 16'hDA81;
reg [15:00] reg_datpt_119 = 16'hB0FB;
reg [15:00] reg_datpt_120 = 16'h7FFF;
reg [15:00] reg_datpt_121 = 16'h4F03;
reg [15:00] reg_datpt_122 = 16'h257D;
reg [15:00] reg_datpt_123 = 16'h09BE;
reg [15:00] reg_datpt_124 = 16'h0000;
reg [15:00] reg_datpt_125 = 16'h09BE;
reg [15:00] reg_datpt_126 = 16'h257D;
reg [15:00] reg_datpt_127 = 16'h4F03;
reg [15:00] reg_datpt_128 = 16'h7FFF;
reg [15:00] reg_datpt_129 = 16'hB0FB;
reg [15:00] reg_datpt_130 = 16'hDA81;
reg [15:00] reg_datpt_131 = 16'hF640;
reg [15:00] reg_datpt_132 = 16'hFFFF;
reg [15:00] reg_datpt_133 = 16'hF640;
reg [15:00] reg_datpt_134 = 16'hDA81;
reg [15:00] reg_datpt_135 = 16'hB0FB;
reg [15:00] reg_datpt_136 = 16'h7FFF;
reg [15:00] reg_datpt_137 = 16'h4F03;
reg [15:00] reg_datpt_138 = 16'h257D;
reg [15:00] reg_datpt_139 = 16'h09BE;
reg [15:00] reg_datpt_140 = 16'h0000;
reg [15:00] reg_datpt_141 = 16'h09BE;
reg [15:00] reg_datpt_142 = 16'h257D;
reg [15:00] reg_datpt_143 = 16'h4F03;
reg [15:00] reg_datpt_144 = 16'h7FFF;
reg [15:00] reg_datpt_145 = 16'hB0FB;
reg [15:00] reg_datpt_146 = 16'hDA81;
reg [15:00] reg_datpt_147 = 16'hF640;
reg [15:00] reg_datpt_148 = 16'hFFFF;
reg [15:00] reg_datpt_149 = 16'hF640;
reg [15:00] reg_datpt_150 = 16'hDA81;
reg [15:00] reg_datpt_151 = 16'hB0FB;
reg [15:00] reg_datpt_152 = 16'h7FFF;
reg [15:00] reg_datpt_153 = 16'h4F03;
reg [15:00] reg_datpt_154 = 16'h257D;
reg [15:00] reg_datpt_155 = 16'h09BE;
reg [15:00] reg_datpt_156 = 16'h0000;
reg [15:00] reg_datpt_157 = 16'h09BE;
reg [15:00] reg_datpt_158 = 16'h257D;
reg [15:00] reg_datpt_159 = 16'h4F03;
reg [15:00] reg_datpt_160 = 16'h7FFF;
reg [15:00] reg_datpt_161 = 16'hB0FB;
reg [15:00] reg_datpt_162 = 16'hDA81;
reg [15:00] reg_datpt_163 = 16'hF640;
reg [15:00] reg_datpt_164 = 16'hFFFF;
reg [15:00] reg_datpt_165 = 16'hF640;
reg [15:00] reg_datpt_166 = 16'hDA81;
reg [15:00] reg_datpt_167 = 16'hB0FB;
reg [15:00] reg_datpt_168 = 16'h7FFF;
reg [15:00] reg_datpt_169 = 16'h4F03;
reg [15:00] reg_datpt_170 = 16'h257D;
reg [15:00] reg_datpt_171 = 16'h09BE;
reg [15:00] reg_datpt_172 = 16'h0000;
reg [15:00] reg_datpt_173 = 16'h09BE;
reg [15:00] reg_datpt_174 = 16'h257D;
reg [15:00] reg_datpt_175 = 16'h4F03;
reg [15:00] reg_datpt_176 = 16'h7FFF;
reg [15:00] reg_datpt_177 = 16'hB0FB;
reg [15:00] reg_datpt_178 = 16'hDA81;
reg [15:00] reg_datpt_179 = 16'hF640;
reg [15:00] reg_datpt_180 = 16'hFFFF;
reg [15:00] reg_datpt_181 = 16'hF640;
reg [15:00] reg_datpt_182 = 16'hDA81;
reg [15:00] reg_datpt_183 = 16'hB0FB;
reg [15:00] reg_datpt_184 = 16'h7FFF;
reg [15:00] reg_datpt_185 = 16'h4F03;
reg [15:00] reg_datpt_186 = 16'h257D;
reg [15:00] reg_datpt_187 = 16'h09BE;
reg [15:00] reg_datpt_188 = 16'h0000;
reg [15:00] reg_datpt_189 = 16'h09BE;
reg [15:00] reg_datpt_190 = 16'h257D;
reg [15:00] reg_datpt_191 = 16'h4F03;
reg [15:00] reg_datpt_192 = 16'h7FFF;
reg [15:00] reg_datpt_193 = 16'hB0FB;
reg [15:00] reg_datpt_194 = 16'hDA81;
reg [15:00] reg_datpt_195 = 16'hF640;
reg [15:00] reg_datpt_196 = 16'hFFFF;
reg [15:00] reg_datpt_197 = 16'hF640;
reg [15:00] reg_datpt_198 = 16'hDA81;
reg [15:00] reg_datpt_199 = 16'hB0FB;
reg [15:00] reg_datpt_200 = 16'h7FFF;
reg [15:00] reg_datpt_201 = 16'h4F03;
reg [15:00] reg_datpt_202 = 16'h257D;
reg [15:00] reg_datpt_203 = 16'h09BE;
reg [15:00] reg_datpt_204 = 16'h0000;
reg [15:00] reg_datpt_205 = 16'h09BE;
reg [15:00] reg_datpt_206 = 16'h257D;
reg [15:00] reg_datpt_207 = 16'h4F03;
reg [15:00] reg_datpt_208 = 16'h7FFF;
reg [15:00] reg_datpt_209 = 16'hB0FB;
reg [15:00] reg_datpt_210 = 16'hDA81;
reg [15:00] reg_datpt_211 = 16'hF640;
reg [15:00] reg_datpt_212 = 16'hFFFF;
reg [15:00] reg_datpt_213 = 16'hF640;
reg [15:00] reg_datpt_214 = 16'hDA81;
reg [15:00] reg_datpt_215 = 16'hB0FB;
reg [15:00] reg_datpt_216 = 16'h7FFF;
reg [15:00] reg_datpt_217 = 16'h4F03;
reg [15:00] reg_datpt_218 = 16'h257D;
reg [15:00] reg_datpt_219 = 16'h09BE;
reg [15:00] reg_datpt_220 = 16'h0000;
reg [15:00] reg_datpt_221 = 16'h09BE;
reg [15:00] reg_datpt_222 = 16'h257D;
reg [15:00] reg_datpt_223 = 16'h4F03;
reg [15:00] reg_datpt_224 = 16'h7FFF;
reg [15:00] reg_datpt_225 = 16'hB0FB;
reg [15:00] reg_datpt_226 = 16'hDA81;
reg [15:00] reg_datpt_227 = 16'hF640;
reg [15:00] reg_datpt_228 = 16'hFFFF;
reg [15:00] reg_datpt_229 = 16'hF640;
reg [15:00] reg_datpt_230 = 16'hDA81;
reg [15:00] reg_datpt_231 = 16'hB0FB;
reg [15:00] reg_datpt_232 = 16'h7FFF;
reg [15:00] reg_datpt_233 = 16'h4F03;
reg [15:00] reg_datpt_234 = 16'h257D;
reg [15:00] reg_datpt_235 = 16'h09BE;
reg [15:00] reg_datpt_236 = 16'h0000;
reg [15:00] reg_datpt_237 = 16'h09BE;
reg [15:00] reg_datpt_238 = 16'h257D;
reg [15:00] reg_datpt_239 = 16'h4F03;
reg [15:00] reg_datpt_240 = 16'h7FFF;
reg [15:00] reg_datpt_241 = 16'hB0FB;
reg [15:00] reg_datpt_242 = 16'hDA81;
reg [15:00] reg_datpt_243 = 16'hF640;
reg [15:00] reg_datpt_244 = 16'hFFFF;
reg [15:00] reg_datpt_245 = 16'hF640;
reg [15:00] reg_datpt_246 = 16'hDA81;
reg [15:00] reg_datpt_247 = 16'hB0FB;
reg [15:00] reg_datpt_248 = 16'h7FFF;
reg [15:00] reg_datpt_249 = 16'h4F03;
reg [15:00] reg_datpt_250 = 16'h257D;
reg [15:00] reg_datpt_251 = 16'h09BE;
reg [15:00] reg_datpt_252 = 16'h0000;
reg [15:00] reg_datpt_253 = 16'h09BE;
reg [15:00] reg_datpt_254 = 16'h257D;
reg [15:00] reg_datpt_255 = 16'h4F03;

reg [7:0] count_i = 8'h0;

always @(posedge CLK or negedge RST)
begin
    if(!RST)                        // Active Low Reset
    begin
        data_pt <= 16'h0;
    end 
    else                            // Reset is High
    begin	                       
        if(Bit == 1'b1)             // Bit-1
        begin 
            case (count_i)
              000 : data_pt <= reg_datpt_000;
              001 : data_pt <= reg_datpt_001;
              002 : data_pt <= reg_datpt_002;
              003 : data_pt <= reg_datpt_003;
              004 : data_pt <= reg_datpt_004;
              005 : data_pt <= reg_datpt_005;
              006 : data_pt <= reg_datpt_006;
              007 : data_pt <= reg_datpt_007;
              008 : data_pt <= reg_datpt_008;
              009 : data_pt <= reg_datpt_009;
              010 : data_pt <= reg_datpt_010;
              011 : data_pt <= reg_datpt_011;
              012 : data_pt <= reg_datpt_012;
              013 : data_pt <= reg_datpt_013;
              014 : data_pt <= reg_datpt_014;
              015 : data_pt <= reg_datpt_015;
              016 : data_pt <= reg_datpt_016;
              017 : data_pt <= reg_datpt_017;
              018 : data_pt <= reg_datpt_018;
              019 : data_pt <= reg_datpt_019;
              020 : data_pt <= reg_datpt_020;
              021 : data_pt <= reg_datpt_021;
              022 : data_pt <= reg_datpt_022;
              023 : data_pt <= reg_datpt_023;
              024 : data_pt <= reg_datpt_024;
              025 : data_pt <= reg_datpt_025;
              026 : data_pt <= reg_datpt_026;
              027 : data_pt <= reg_datpt_027;
              028 : data_pt <= reg_datpt_028;
              029 : data_pt <= reg_datpt_029;
              030 : data_pt <= reg_datpt_030;
              031 : data_pt <= reg_datpt_031;
              032 : data_pt <= reg_datpt_032;
              033 : data_pt <= reg_datpt_033;
              034 : data_pt <= reg_datpt_034;
              035 : data_pt <= reg_datpt_035;
              036 : data_pt <= reg_datpt_036;
              037 : data_pt <= reg_datpt_037;
              038 : data_pt <= reg_datpt_038;
              039 : data_pt <= reg_datpt_039;
              040 : data_pt <= reg_datpt_040;
              041 : data_pt <= reg_datpt_041;
              042 : data_pt <= reg_datpt_042;
              043 : data_pt <= reg_datpt_043;
              044 : data_pt <= reg_datpt_044;
              045 : data_pt <= reg_datpt_045;
              046 : data_pt <= reg_datpt_046;
              047 : data_pt <= reg_datpt_047;
              048 : data_pt <= reg_datpt_048;
              049 : data_pt <= reg_datpt_049;
              050 : data_pt <= reg_datpt_050;
              051 : data_pt <= reg_datpt_051;
              052 : data_pt <= reg_datpt_052;
              053 : data_pt <= reg_datpt_053;
              054 : data_pt <= reg_datpt_054;
              055 : data_pt <= reg_datpt_055;
              056 : data_pt <= reg_datpt_056;
              057 : data_pt <= reg_datpt_057;
              058 : data_pt <= reg_datpt_058;
              059 : data_pt <= reg_datpt_059;
              060 : data_pt <= reg_datpt_060;
              061 : data_pt <= reg_datpt_061;
              062 : data_pt <= reg_datpt_062;
              063 : data_pt <= reg_datpt_063;
              064 : data_pt <= reg_datpt_064;
              065 : data_pt <= reg_datpt_065;
              066 : data_pt <= reg_datpt_066;
              067 : data_pt <= reg_datpt_067;
              068 : data_pt <= reg_datpt_068;
              069 : data_pt <= reg_datpt_069;
              070 : data_pt <= reg_datpt_070;
              071 : data_pt <= reg_datpt_071;
              072 : data_pt <= reg_datpt_072;
              073 : data_pt <= reg_datpt_073;
              074 : data_pt <= reg_datpt_074;
              075 : data_pt <= reg_datpt_075;
              076 : data_pt <= reg_datpt_076;
              077 : data_pt <= reg_datpt_077;
              078 : data_pt <= reg_datpt_078;
              079 : data_pt <= reg_datpt_079;
              080 : data_pt <= reg_datpt_080;
              081 : data_pt <= reg_datpt_081;
              082 : data_pt <= reg_datpt_082;
              083 : data_pt <= reg_datpt_083;
              084 : data_pt <= reg_datpt_084;
              085 : data_pt <= reg_datpt_085;
              086 : data_pt <= reg_datpt_086;
              087 : data_pt <= reg_datpt_087;
              088 : data_pt <= reg_datpt_088;
              089 : data_pt <= reg_datpt_089;
              090 : data_pt <= reg_datpt_090;
              091 : data_pt <= reg_datpt_091;
              092 : data_pt <= reg_datpt_092;
              093 : data_pt <= reg_datpt_093;
              094 : data_pt <= reg_datpt_094;
              095 : data_pt <= reg_datpt_095;
              096 : data_pt <= reg_datpt_096;
              097 : data_pt <= reg_datpt_097;
              098 : data_pt <= reg_datpt_098;
              099 : data_pt <= reg_datpt_099;
              100 : data_pt <= reg_datpt_100;
              101 : data_pt <= reg_datpt_101;
              102 : data_pt <= reg_datpt_102;
              103 : data_pt <= reg_datpt_103;
              104 : data_pt <= reg_datpt_104;
              105 : data_pt <= reg_datpt_105;
              106 : data_pt <= reg_datpt_106;
              107 : data_pt <= reg_datpt_107;
              108 : data_pt <= reg_datpt_108;
              109 : data_pt <= reg_datpt_109;
              110 : data_pt <= reg_datpt_110;
              111 : data_pt <= reg_datpt_111;
              112 : data_pt <= reg_datpt_112;
              113 : data_pt <= reg_datpt_113;
              114 : data_pt <= reg_datpt_114;
              115 : data_pt <= reg_datpt_115;
              116 : data_pt <= reg_datpt_116;
              117 : data_pt <= reg_datpt_117;
              118 : data_pt <= reg_datpt_118;
              119 : data_pt <= reg_datpt_119;
              120 : data_pt <= reg_datpt_120;
              121 : data_pt <= reg_datpt_121;
              122 : data_pt <= reg_datpt_122;
              123 : data_pt <= reg_datpt_123;
              124 : data_pt <= reg_datpt_124;
              125 : data_pt <= reg_datpt_125;
              126 : data_pt <= reg_datpt_126;
              127 : data_pt <= reg_datpt_127;
              128 : data_pt <= reg_datpt_128;
              129 : data_pt <= reg_datpt_129;
              130 : data_pt <= reg_datpt_130;
              131 : data_pt <= reg_datpt_131;
              132 : data_pt <= reg_datpt_132;
              133 : data_pt <= reg_datpt_133;
              134 : data_pt <= reg_datpt_134;
              135 : data_pt <= reg_datpt_135;
              136 : data_pt <= reg_datpt_136;
              137 : data_pt <= reg_datpt_137;
              138 : data_pt <= reg_datpt_138;
              139 : data_pt <= reg_datpt_139;
              140 : data_pt <= reg_datpt_140;
              141 : data_pt <= reg_datpt_141;
              142 : data_pt <= reg_datpt_142;
              143 : data_pt <= reg_datpt_143;
              144 : data_pt <= reg_datpt_144;
              145 : data_pt <= reg_datpt_145;
              146 : data_pt <= reg_datpt_146;
              147 : data_pt <= reg_datpt_147;
              148 : data_pt <= reg_datpt_148;
              149 : data_pt <= reg_datpt_149;
              150 : data_pt <= reg_datpt_150;
              151 : data_pt <= reg_datpt_151;
              152 : data_pt <= reg_datpt_152;
              153 : data_pt <= reg_datpt_153;
              154 : data_pt <= reg_datpt_154;
              155 : data_pt <= reg_datpt_155;
              156 : data_pt <= reg_datpt_156;
              157 : data_pt <= reg_datpt_157;
              158 : data_pt <= reg_datpt_158;
              159 : data_pt <= reg_datpt_159;
              160 : data_pt <= reg_datpt_160;
              161 : data_pt <= reg_datpt_161;
              162 : data_pt <= reg_datpt_162;
              163 : data_pt <= reg_datpt_163;
              164 : data_pt <= reg_datpt_164;
              165 : data_pt <= reg_datpt_165;
              166 : data_pt <= reg_datpt_166;
              167 : data_pt <= reg_datpt_167;
              168 : data_pt <= reg_datpt_168;
              169 : data_pt <= reg_datpt_169;
              170 : data_pt <= reg_datpt_170;
              171 : data_pt <= reg_datpt_171;
              172 : data_pt <= reg_datpt_172;
              173 : data_pt <= reg_datpt_173;
              174 : data_pt <= reg_datpt_174;
              175 : data_pt <= reg_datpt_175;
              176 : data_pt <= reg_datpt_176;
              177 : data_pt <= reg_datpt_177;
              178 : data_pt <= reg_datpt_178;
              179 : data_pt <= reg_datpt_179;
              180 : data_pt <= reg_datpt_180;
              181 : data_pt <= reg_datpt_181;
              182 : data_pt <= reg_datpt_182;
              183 : data_pt <= reg_datpt_183;
              184 : data_pt <= reg_datpt_184;
              185 : data_pt <= reg_datpt_185;
              186 : data_pt <= reg_datpt_186;
              187 : data_pt <= reg_datpt_187;
              188 : data_pt <= reg_datpt_188;
              189 : data_pt <= reg_datpt_189;
              190 : data_pt <= reg_datpt_190;
              191 : data_pt <= reg_datpt_191;
              192 : data_pt <= reg_datpt_192;
              193 : data_pt <= reg_datpt_193;
              194 : data_pt <= reg_datpt_194;
              195 : data_pt <= reg_datpt_195;
              196 : data_pt <= reg_datpt_196;
              197 : data_pt <= reg_datpt_197;
              198 : data_pt <= reg_datpt_198;
              199 : data_pt <= reg_datpt_199;
              200 : data_pt <= reg_datpt_200;
              201 : data_pt <= reg_datpt_201;
              202 : data_pt <= reg_datpt_202;
              203 : data_pt <= reg_datpt_203;
              204 : data_pt <= reg_datpt_204;
              205 : data_pt <= reg_datpt_205;
              206 : data_pt <= reg_datpt_206;
              207 : data_pt <= reg_datpt_207;
              208 : data_pt <= reg_datpt_208;
              209 : data_pt <= reg_datpt_209;
              210 : data_pt <= reg_datpt_210;
              211 : data_pt <= reg_datpt_211;
              212 : data_pt <= reg_datpt_212;
              213 : data_pt <= reg_datpt_213;
              214 : data_pt <= reg_datpt_214;
              215 : data_pt <= reg_datpt_215;
              216 : data_pt <= reg_datpt_216;
              217 : data_pt <= reg_datpt_217;
              218 : data_pt <= reg_datpt_218;
              219 : data_pt <= reg_datpt_219;
              220 : data_pt <= reg_datpt_220;
              221 : data_pt <= reg_datpt_221;
              222 : data_pt <= reg_datpt_222;
              223 : data_pt <= reg_datpt_223;
              224 : data_pt <= reg_datpt_224;
              225 : data_pt <= reg_datpt_225;
              226 : data_pt <= reg_datpt_226;
              227 : data_pt <= reg_datpt_227;
              228 : data_pt <= reg_datpt_228;
              229 : data_pt <= reg_datpt_229;
              230 : data_pt <= reg_datpt_230;
              231 : data_pt <= reg_datpt_231;
              232 : data_pt <= reg_datpt_232;
              233 : data_pt <= reg_datpt_233;
              234 : data_pt <= reg_datpt_234;
              235 : data_pt <= reg_datpt_235;
              236 : data_pt <= reg_datpt_236;
              237 : data_pt <= reg_datpt_237;
              238 : data_pt <= reg_datpt_238;
              239 : data_pt <= reg_datpt_239;
              240 : data_pt <= reg_datpt_240;
              241 : data_pt <= reg_datpt_241;
              242 : data_pt <= reg_datpt_242;
              243 : data_pt <= reg_datpt_243;
              244 : data_pt <= reg_datpt_244;
              245 : data_pt <= reg_datpt_245;
              246 : data_pt <= reg_datpt_246;
              247 : data_pt <= reg_datpt_247;
              248 : data_pt <= reg_datpt_248;
              249 : data_pt <= reg_datpt_249;
              250 : data_pt <= reg_datpt_250;
              251 : data_pt <= reg_datpt_251;
              252 : data_pt <= reg_datpt_252;
              253 : data_pt <= reg_datpt_253;
              254 : data_pt <= reg_datpt_254;
              255 : data_pt <= reg_datpt_255;
            endcase
        end     
        else if(Bit == 1'b0)
        begin
            case (count_i)      // Bit-0, Divide Amplitude by 2
              000 : data_pt <= reg_datpt_000 >> 1;
              001 : data_pt <= reg_datpt_001 >> 1;
              002 : data_pt <= reg_datpt_002 >> 1;
              003 : data_pt <= reg_datpt_003 >> 1;
              004 : data_pt <= reg_datpt_004 >> 1;
              005 : data_pt <= reg_datpt_005 >> 1;
              006 : data_pt <= reg_datpt_006 >> 1;
              007 : data_pt <= reg_datpt_007 >> 1;
              008 : data_pt <= reg_datpt_008 >> 1;
              009 : data_pt <= reg_datpt_009 >> 1;
              010 : data_pt <= reg_datpt_010 >> 1;
              011 : data_pt <= reg_datpt_011 >> 1;
              012 : data_pt <= reg_datpt_012 >> 1;
              013 : data_pt <= reg_datpt_013 >> 1;
              014 : data_pt <= reg_datpt_014 >> 1;
              015 : data_pt <= reg_datpt_015 >> 1;
              016 : data_pt <= reg_datpt_016 >> 1;
              017 : data_pt <= reg_datpt_017 >> 1;
              018 : data_pt <= reg_datpt_018 >> 1;
              019 : data_pt <= reg_datpt_019 >> 1;
              020 : data_pt <= reg_datpt_020 >> 1;
              021 : data_pt <= reg_datpt_021 >> 1;
              022 : data_pt <= reg_datpt_022 >> 1;
              023 : data_pt <= reg_datpt_023 >> 1;
              024 : data_pt <= reg_datpt_024 >> 1;
              025 : data_pt <= reg_datpt_025 >> 1;
              026 : data_pt <= reg_datpt_026 >> 1;
              027 : data_pt <= reg_datpt_027 >> 1;
              028 : data_pt <= reg_datpt_028 >> 1;
              029 : data_pt <= reg_datpt_029 >> 1;
              030 : data_pt <= reg_datpt_030 >> 1;
              031 : data_pt <= reg_datpt_031 >> 1;
              032 : data_pt <= reg_datpt_032 >> 1;
              033 : data_pt <= reg_datpt_033 >> 1;
              034 : data_pt <= reg_datpt_034 >> 1;
              035 : data_pt <= reg_datpt_035 >> 1;
              036 : data_pt <= reg_datpt_036 >> 1;
              037 : data_pt <= reg_datpt_037 >> 1;
              038 : data_pt <= reg_datpt_038 >> 1;
              039 : data_pt <= reg_datpt_039 >> 1;
              040 : data_pt <= reg_datpt_040 >> 1;
              041 : data_pt <= reg_datpt_041 >> 1;
              042 : data_pt <= reg_datpt_042 >> 1;
              043 : data_pt <= reg_datpt_043 >> 1;
              044 : data_pt <= reg_datpt_044 >> 1;
              045 : data_pt <= reg_datpt_045 >> 1;
              046 : data_pt <= reg_datpt_046 >> 1;
              047 : data_pt <= reg_datpt_047 >> 1;
              048 : data_pt <= reg_datpt_048 >> 1;
              049 : data_pt <= reg_datpt_049 >> 1;
              050 : data_pt <= reg_datpt_050 >> 1;
              051 : data_pt <= reg_datpt_051 >> 1;
              052 : data_pt <= reg_datpt_052 >> 1;
              053 : data_pt <= reg_datpt_053 >> 1;
              054 : data_pt <= reg_datpt_054 >> 1;
              055 : data_pt <= reg_datpt_055 >> 1;
              056 : data_pt <= reg_datpt_056 >> 1;
              057 : data_pt <= reg_datpt_057 >> 1;
              058 : data_pt <= reg_datpt_058 >> 1;
              059 : data_pt <= reg_datpt_059 >> 1;
              060 : data_pt <= reg_datpt_060 >> 1;
              061 : data_pt <= reg_datpt_061 >> 1;
              062 : data_pt <= reg_datpt_062 >> 1;
              063 : data_pt <= reg_datpt_063 >> 1;
              064 : data_pt <= reg_datpt_064 >> 1;
              065 : data_pt <= reg_datpt_065 >> 1;
              066 : data_pt <= reg_datpt_066 >> 1;
              067 : data_pt <= reg_datpt_067 >> 1;
              068 : data_pt <= reg_datpt_068 >> 1;
              069 : data_pt <= reg_datpt_069 >> 1;
              070 : data_pt <= reg_datpt_070 >> 1;
              071 : data_pt <= reg_datpt_071 >> 1;
              072 : data_pt <= reg_datpt_072 >> 1;
              073 : data_pt <= reg_datpt_073 >> 1;
              074 : data_pt <= reg_datpt_074 >> 1;
              075 : data_pt <= reg_datpt_075 >> 1;
              076 : data_pt <= reg_datpt_076 >> 1;
              077 : data_pt <= reg_datpt_077 >> 1;
              078 : data_pt <= reg_datpt_078 >> 1;
              079 : data_pt <= reg_datpt_079 >> 1;
              080 : data_pt <= reg_datpt_080 >> 1;
              081 : data_pt <= reg_datpt_081 >> 1;
              082 : data_pt <= reg_datpt_082 >> 1;
              083 : data_pt <= reg_datpt_083 >> 1;
              084 : data_pt <= reg_datpt_084 >> 1;
              085 : data_pt <= reg_datpt_085 >> 1;
              086 : data_pt <= reg_datpt_086 >> 1;
              087 : data_pt <= reg_datpt_087 >> 1;
              088 : data_pt <= reg_datpt_088 >> 1;
              089 : data_pt <= reg_datpt_089 >> 1;
              090 : data_pt <= reg_datpt_090 >> 1;
              091 : data_pt <= reg_datpt_091 >> 1;
              092 : data_pt <= reg_datpt_092 >> 1;
              093 : data_pt <= reg_datpt_093 >> 1;
              094 : data_pt <= reg_datpt_094 >> 1;
              095 : data_pt <= reg_datpt_095 >> 1;
              096 : data_pt <= reg_datpt_096 >> 1;
              097 : data_pt <= reg_datpt_097 >> 1;
              098 : data_pt <= reg_datpt_098 >> 1;
              099 : data_pt <= reg_datpt_099 >> 1;
              100 : data_pt <= reg_datpt_100 >> 1;
              101 : data_pt <= reg_datpt_101 >> 1;
              102 : data_pt <= reg_datpt_102 >> 1;
              103 : data_pt <= reg_datpt_103 >> 1;
              104 : data_pt <= reg_datpt_104 >> 1;
              105 : data_pt <= reg_datpt_105 >> 1;
              106 : data_pt <= reg_datpt_106 >> 1;
              107 : data_pt <= reg_datpt_107 >> 1;
              108 : data_pt <= reg_datpt_108 >> 1;
              109 : data_pt <= reg_datpt_109 >> 1;
              110 : data_pt <= reg_datpt_110 >> 1;
              111 : data_pt <= reg_datpt_111 >> 1;
              112 : data_pt <= reg_datpt_112 >> 1;
              113 : data_pt <= reg_datpt_113 >> 1;
              114 : data_pt <= reg_datpt_114 >> 1;
              115 : data_pt <= reg_datpt_115 >> 1;
              116 : data_pt <= reg_datpt_116 >> 1;
              117 : data_pt <= reg_datpt_117 >> 1;
              118 : data_pt <= reg_datpt_118 >> 1;
              119 : data_pt <= reg_datpt_119 >> 1;
              120 : data_pt <= reg_datpt_120 >> 1;
              121 : data_pt <= reg_datpt_121 >> 1;
              122 : data_pt <= reg_datpt_122 >> 1;
              123 : data_pt <= reg_datpt_123 >> 1;
              124 : data_pt <= reg_datpt_124 >> 1;
              125 : data_pt <= reg_datpt_125 >> 1;
              126 : data_pt <= reg_datpt_126 >> 1;
              127 : data_pt <= reg_datpt_127 >> 1;
              128 : data_pt <= reg_datpt_128 >> 1;
              129 : data_pt <= reg_datpt_129 >> 1;
              130 : data_pt <= reg_datpt_130 >> 1;
              131 : data_pt <= reg_datpt_131 >> 1;
              132 : data_pt <= reg_datpt_132 >> 1;
              133 : data_pt <= reg_datpt_133 >> 1;
              134 : data_pt <= reg_datpt_134 >> 1;
              135 : data_pt <= reg_datpt_135 >> 1;
              136 : data_pt <= reg_datpt_136 >> 1;
              137 : data_pt <= reg_datpt_137 >> 1;
              138 : data_pt <= reg_datpt_138 >> 1;
              139 : data_pt <= reg_datpt_139 >> 1;
              140 : data_pt <= reg_datpt_140 >> 1;
              141 : data_pt <= reg_datpt_141 >> 1;
              142 : data_pt <= reg_datpt_142 >> 1;
              143 : data_pt <= reg_datpt_143 >> 1;
              144 : data_pt <= reg_datpt_144 >> 1;
              145 : data_pt <= reg_datpt_145 >> 1;
              146 : data_pt <= reg_datpt_146 >> 1;
              147 : data_pt <= reg_datpt_147 >> 1;
              148 : data_pt <= reg_datpt_148 >> 1;
              149 : data_pt <= reg_datpt_149 >> 1;
              150 : data_pt <= reg_datpt_150 >> 1;
              151 : data_pt <= reg_datpt_151 >> 1;
              152 : data_pt <= reg_datpt_152 >> 1;
              153 : data_pt <= reg_datpt_153 >> 1;
              154 : data_pt <= reg_datpt_154 >> 1;
              155 : data_pt <= reg_datpt_155 >> 1;
              156 : data_pt <= reg_datpt_156 >> 1;
              157 : data_pt <= reg_datpt_157 >> 1;
              158 : data_pt <= reg_datpt_158 >> 1;
              159 : data_pt <= reg_datpt_159 >> 1;
              160 : data_pt <= reg_datpt_160 >> 1;
              161 : data_pt <= reg_datpt_161 >> 1;
              162 : data_pt <= reg_datpt_162 >> 1;
              163 : data_pt <= reg_datpt_163 >> 1;
              164 : data_pt <= reg_datpt_164 >> 1;
              165 : data_pt <= reg_datpt_165 >> 1;
              166 : data_pt <= reg_datpt_166 >> 1;
              167 : data_pt <= reg_datpt_167 >> 1;
              168 : data_pt <= reg_datpt_168 >> 1;
              169 : data_pt <= reg_datpt_169 >> 1;
              170 : data_pt <= reg_datpt_170 >> 1;
              171 : data_pt <= reg_datpt_171 >> 1;
              172 : data_pt <= reg_datpt_172 >> 1;
              173 : data_pt <= reg_datpt_173 >> 1;
              174 : data_pt <= reg_datpt_174 >> 1;
              175 : data_pt <= reg_datpt_175 >> 1;
              176 : data_pt <= reg_datpt_176 >> 1;
              177 : data_pt <= reg_datpt_177 >> 1;
              178 : data_pt <= reg_datpt_178 >> 1;
              179 : data_pt <= reg_datpt_179 >> 1;
              180 : data_pt <= reg_datpt_180 >> 1;
              181 : data_pt <= reg_datpt_181 >> 1;
              182 : data_pt <= reg_datpt_182 >> 1;
              183 : data_pt <= reg_datpt_183 >> 1;
              184 : data_pt <= reg_datpt_184 >> 1;
              185 : data_pt <= reg_datpt_185 >> 1;
              186 : data_pt <= reg_datpt_186 >> 1;
              187 : data_pt <= reg_datpt_187 >> 1;
              188 : data_pt <= reg_datpt_188 >> 1;
              189 : data_pt <= reg_datpt_189 >> 1;
              190 : data_pt <= reg_datpt_190 >> 1;
              191 : data_pt <= reg_datpt_191 >> 1;
              192 : data_pt <= reg_datpt_192 >> 1;
              193 : data_pt <= reg_datpt_193 >> 1;
              194 : data_pt <= reg_datpt_194 >> 1;
              195 : data_pt <= reg_datpt_195 >> 1;
              196 : data_pt <= reg_datpt_196 >> 1;
              197 : data_pt <= reg_datpt_197 >> 1;
              198 : data_pt <= reg_datpt_198 >> 1;
              199 : data_pt <= reg_datpt_199 >> 1;
              200 : data_pt <= reg_datpt_200 >> 1;
              201 : data_pt <= reg_datpt_201 >> 1;
              202 : data_pt <= reg_datpt_202 >> 1;
              203 : data_pt <= reg_datpt_203 >> 1;
              204 : data_pt <= reg_datpt_204 >> 1;
              205 : data_pt <= reg_datpt_205 >> 1;
              206 : data_pt <= reg_datpt_206 >> 1;
              207 : data_pt <= reg_datpt_207 >> 1;
              208 : data_pt <= reg_datpt_208 >> 1;
              209 : data_pt <= reg_datpt_209 >> 1;
              210 : data_pt <= reg_datpt_210 >> 1;
              211 : data_pt <= reg_datpt_211 >> 1;
              212 : data_pt <= reg_datpt_212 >> 1;
              213 : data_pt <= reg_datpt_213 >> 1;
              214 : data_pt <= reg_datpt_214 >> 1;
              215 : data_pt <= reg_datpt_215 >> 1;
              216 : data_pt <= reg_datpt_216 >> 1;
              217 : data_pt <= reg_datpt_217 >> 1;
              218 : data_pt <= reg_datpt_218 >> 1;
              219 : data_pt <= reg_datpt_219 >> 1;
              220 : data_pt <= reg_datpt_220 >> 1;
              221 : data_pt <= reg_datpt_221 >> 1;
              222 : data_pt <= reg_datpt_222 >> 1;
              223 : data_pt <= reg_datpt_223 >> 1;
              224 : data_pt <= reg_datpt_224 >> 1;
              225 : data_pt <= reg_datpt_225 >> 1;
              226 : data_pt <= reg_datpt_226 >> 1;
              227 : data_pt <= reg_datpt_227 >> 1;
              228 : data_pt <= reg_datpt_228 >> 1;
              229 : data_pt <= reg_datpt_229 >> 1;
              230 : data_pt <= reg_datpt_230 >> 1;
              231 : data_pt <= reg_datpt_231 >> 1;
              232 : data_pt <= reg_datpt_232 >> 1;
              233 : data_pt <= reg_datpt_233 >> 1;
              234 : data_pt <= reg_datpt_234 >> 1;
              235 : data_pt <= reg_datpt_235 >> 1;
              236 : data_pt <= reg_datpt_236 >> 1;
              237 : data_pt <= reg_datpt_237 >> 1;
              238 : data_pt <= reg_datpt_238 >> 1;
              239 : data_pt <= reg_datpt_239 >> 1;
              240 : data_pt <= reg_datpt_240 >> 1;
              241 : data_pt <= reg_datpt_241 >> 1;
              242 : data_pt <= reg_datpt_242 >> 1;
              243 : data_pt <= reg_datpt_243 >> 1;
              244 : data_pt <= reg_datpt_244 >> 1;
              245 : data_pt <= reg_datpt_245 >> 1;
              246 : data_pt <= reg_datpt_246 >> 1;
              247 : data_pt <= reg_datpt_247 >> 1;
              248 : data_pt <= reg_datpt_248 >> 1;
              249 : data_pt <= reg_datpt_249 >> 1;
              250 : data_pt <= reg_datpt_250 >> 1;
              251 : data_pt <= reg_datpt_251 >> 1;
              252 : data_pt <= reg_datpt_252 >> 1;
              253 : data_pt <= reg_datpt_253 >> 1;
              254 : data_pt <= reg_datpt_254 >> 1;
              255 : data_pt <= reg_datpt_255 >> 1;
            endcase         
        end
        count_i <= count_i + 8'h1;  
    end
    if(count_i == 255)
        dFLAG <= 1'b1;
    else
        dFLAG <= 1'b0;
end
endmodule
